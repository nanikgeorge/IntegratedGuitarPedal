* NGSPICE file created from sbi_flat.ext - technology: sky130A

.subckt test_inverter IN OUT VSS VDD
X0 IN OUT VSS sky130_fd_pr__res_xhigh_po_0p35 l=26.11
X1 OUT.t0 IN.t1 VSS.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X2 IN OUT VSS.t2 sky130_fd_pr__res_xhigh_po_0p35 l=0.16
X3 OUT.t1 IN.t2 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
R0 IN.n0 IN.t2 120.174
R1 IN.n1 IN.t1 118.005
R2 IN.n2 IN 0.455045
R3 IN.n0 IN 0.229416
R4 IN.n2 IN.n1 0.0745741
R5 IN IN.n2 0.0174753
R6 IN.n1 IN.n0 0.0128457
R7 OUT.n0 OUT.t1 228.32
R8 OUT OUT.t0 83.7895
R9 OUT.n1 OUT.n0 0.417167
R10 OUT.n0 OUT 0.354667
R11 OUT OUT.n1 0.292167
R12 OUT.n1 OUT 0.0272857
R13 VSS.n1 VSS.n0 250.325
R14 VSS.n1 VSS.t1 84.039
R15 VSS.n0 VSS.t2 50.0542
R16 VSS.n0 VSS.t0 20.7127
R17 VSS VSS.n1 0.2005
R18 VDD.n0 VDD.t0 658.12
R19 VDD.n0 VDD.t1 228.59
R20 VDD VDD.n0 0.163
C0 OUT VDD 0.119038f
C1 OUT IN 0.156189f
C2 VDD IN 0.330567f
C3 OUT VSS 1.01935f
C4 IN VSS 1.54313f
C5 VDD VSS 0.96518f
.ends

