magic
tech sky130A
magscale 1 2
timestamp 1713408040
<< locali >>
rect -50 1000 800 1050
rect -50 600 20 1000
rect 720 880 800 1000
rect 80 680 150 850
rect 600 680 660 850
rect 80 600 280 680
rect 220 520 280 600
rect 460 600 660 680
rect 720 840 1000 880
rect 720 660 880 840
rect 980 660 1000 840
rect 720 620 1000 660
rect 460 520 520 600
rect 220 440 520 520
rect -50 20 20 400
rect 80 200 150 400
rect 320 160 420 440
rect 600 200 660 400
rect 720 360 1000 400
rect 720 180 880 360
rect 980 180 1000 360
rect 720 140 1000 180
rect 720 20 800 140
rect -50 -50 800 20
<< viali >>
rect 880 660 980 840
rect 880 180 980 360
<< metal1 >>
rect 140 1180 600 1200
rect 140 1000 160 1180
rect 580 1000 600 1180
rect 140 900 600 1000
rect -80 840 180 860
rect -80 660 -60 840
rect 160 660 180 840
rect -80 640 180 660
rect 320 560 420 860
rect 560 840 820 860
rect 560 660 580 840
rect 800 660 820 840
rect 560 640 820 660
rect 860 840 1300 860
rect 860 660 880 840
rect 980 660 1300 840
rect 860 640 1300 660
rect 60 480 680 560
rect 60 380 160 480
rect 580 380 680 480
rect -80 360 180 380
rect -80 180 -60 360
rect 160 180 180 360
rect -80 160 180 180
rect 560 360 820 380
rect 560 180 580 360
rect 800 180 820 360
rect 560 160 820 180
rect 860 360 1300 380
rect 860 180 880 360
rect 980 180 1300 360
rect 860 160 1300 180
rect 140 20 600 120
rect 140 -160 160 20
rect 580 -160 600 20
rect 140 -180 600 -160
<< via1 >>
rect 160 1000 580 1180
rect -60 660 160 840
rect 580 660 800 840
rect -60 180 160 360
rect 580 180 800 360
rect 160 -160 580 20
<< metal2 >>
rect -380 1180 1000 1200
rect -380 1000 160 1180
rect 580 1000 1000 1180
rect -380 980 1000 1000
rect -380 840 1000 860
rect -380 660 -60 840
rect 160 660 580 840
rect 800 660 1000 840
rect -380 640 1000 660
rect -380 360 1000 380
rect -380 180 -60 360
rect 160 180 580 360
rect 800 180 1000 360
rect -380 160 1000 180
rect -380 20 1000 40
rect -380 -160 160 20
rect 580 -160 1000 20
rect -380 -180 1000 -160
use sky130_fd_pr__nfet_01v8_7HRXTK  sky130_fd_pr__nfet_01v8_7HRXTK_0
timestamp 1713395545
transform 1 0 372 0 1 226
box -425 -279 425 279
use sky130_fd_pr__pfet_01v8_UNVJW6  sky130_fd_pr__pfet_01v8_UNVJW6_0
timestamp 1713395545
transform 1 0 372 0 1 789
box -425 -284 425 284
<< labels >>
flabel metal2 -380 640 -60 860 0 FreeSans 1600 0 0 0 IN
port 1 nsew
flabel metal2 -380 160 -60 380 0 FreeSans 1600 0 0 0 OUT
port 2 nsew
flabel metal2 -380 980 160 1200 0 FreeSans 1600 0 0 0 CTRLB
port 4 nsew
flabel metal2 -380 -180 160 40 0 FreeSans 1600 0 0 0 CTRL
port 3 nsew
flabel metal1 980 640 1300 860 0 FreeSans 1600 0 0 0 VDD
flabel metal1 980 160 1300 380 0 FreeSans 1600 0 0 0 VSS
<< end >>
