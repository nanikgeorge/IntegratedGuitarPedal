magic
tech sky130A
magscale 1 2
timestamp 1713223699
<< nmos >>
rect -745 -19 -545 81
rect -487 -19 -287 81
rect -229 -19 -29 81
rect 29 -19 229 81
rect 287 -19 487 81
rect 545 -19 745 81
<< ndiff >>
rect -803 69 -745 81
rect -803 -7 -791 69
rect -757 -7 -745 69
rect -803 -19 -745 -7
rect -545 69 -487 81
rect -545 -7 -533 69
rect -499 -7 -487 69
rect -545 -19 -487 -7
rect -287 69 -229 81
rect -287 -7 -275 69
rect -241 -7 -229 69
rect -287 -19 -229 -7
rect -29 69 29 81
rect -29 -7 -17 69
rect 17 -7 29 69
rect -29 -19 29 -7
rect 229 69 287 81
rect 229 -7 241 69
rect 275 -7 287 69
rect 229 -19 287 -7
rect 487 69 545 81
rect 487 -7 499 69
rect 533 -7 545 69
rect 487 -19 545 -7
rect 745 69 803 81
rect 745 -7 757 69
rect 791 -7 803 69
rect 745 -19 803 -7
<< ndiffc >>
rect -791 -7 -757 69
rect -533 -7 -499 69
rect -275 -7 -241 69
rect -17 -7 17 69
rect 241 -7 275 69
rect 499 -7 533 69
rect 757 -7 791 69
<< poly >>
rect -745 81 -545 107
rect -487 81 -287 107
rect -229 81 -29 107
rect 29 81 229 107
rect 287 81 487 107
rect 545 81 745 107
rect -745 -57 -545 -19
rect -745 -91 -729 -57
rect -561 -91 -545 -57
rect -745 -107 -545 -91
rect -487 -57 -287 -19
rect -487 -91 -471 -57
rect -303 -91 -287 -57
rect -487 -107 -287 -91
rect -229 -57 -29 -19
rect -229 -91 -213 -57
rect -45 -91 -29 -57
rect -229 -107 -29 -91
rect 29 -57 229 -19
rect 29 -91 45 -57
rect 213 -91 229 -57
rect 29 -107 229 -91
rect 287 -57 487 -19
rect 287 -91 303 -57
rect 471 -91 487 -57
rect 287 -107 487 -91
rect 545 -57 745 -19
rect 545 -91 561 -57
rect 729 -91 745 -57
rect 545 -107 745 -91
<< polycont >>
rect -729 -91 -561 -57
rect -471 -91 -303 -57
rect -213 -91 -45 -57
rect 45 -91 213 -57
rect 303 -91 471 -57
rect 561 -91 729 -57
<< locali >>
rect -791 69 -757 85
rect -791 -23 -757 -7
rect -533 69 -499 85
rect -533 -23 -499 -7
rect -275 69 -241 85
rect -275 -23 -241 -7
rect -17 69 17 85
rect -17 -23 17 -7
rect 241 69 275 85
rect 241 -23 275 -7
rect 499 69 533 85
rect 499 -23 533 -7
rect 757 69 791 85
rect 757 -23 791 -7
rect -745 -91 -729 -57
rect -561 -91 -545 -57
rect -487 -91 -471 -57
rect -303 -91 -287 -57
rect -229 -91 -213 -57
rect -45 -91 -29 -57
rect 29 -91 45 -57
rect 213 -91 229 -57
rect 287 -91 303 -57
rect 471 -91 487 -57
rect 545 -91 561 -57
rect 729 -91 745 -57
<< viali >>
rect -791 -7 -757 69
rect -533 -7 -499 69
rect -275 -7 -241 69
rect -17 -7 17 69
rect 241 -7 275 69
rect 499 -7 533 69
rect 757 -7 791 69
rect -729 -91 -561 -57
rect -471 -91 -303 -57
rect -213 -91 -45 -57
rect 45 -91 213 -57
rect 303 -91 471 -57
rect 561 -91 729 -57
<< metal1 >>
rect -797 69 -751 81
rect -797 -7 -791 69
rect -757 -7 -751 69
rect -797 -19 -751 -7
rect -539 69 -493 81
rect -539 -7 -533 69
rect -499 -7 -493 69
rect -539 -19 -493 -7
rect -281 69 -235 81
rect -281 -7 -275 69
rect -241 -7 -235 69
rect -281 -19 -235 -7
rect -23 69 23 81
rect -23 -7 -17 69
rect 17 -7 23 69
rect -23 -19 23 -7
rect 235 69 281 81
rect 235 -7 241 69
rect 275 -7 281 69
rect 235 -19 281 -7
rect 493 69 539 81
rect 493 -7 499 69
rect 533 -7 539 69
rect 493 -19 539 -7
rect 751 69 797 81
rect 751 -7 757 69
rect 791 -7 797 69
rect 751 -19 797 -7
rect -741 -57 -549 -51
rect -741 -91 -729 -57
rect -561 -91 -549 -57
rect -741 -97 -549 -91
rect -483 -57 -291 -51
rect -483 -91 -471 -57
rect -303 -91 -291 -57
rect -483 -97 -291 -91
rect -225 -57 -33 -51
rect -225 -91 -213 -57
rect -45 -91 -33 -57
rect -225 -97 -33 -91
rect 33 -57 225 -51
rect 33 -91 45 -57
rect 213 -91 225 -57
rect 33 -97 225 -91
rect 291 -57 483 -51
rect 291 -91 303 -57
rect 471 -91 483 -57
rect 291 -97 483 -91
rect 549 -57 741 -51
rect 549 -91 561 -57
rect 729 -91 741 -57
rect 549 -97 741 -91
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.5 l 1 m 1 nf 6 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
