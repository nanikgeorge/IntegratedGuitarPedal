magic
tech sky130A
magscale 1 2
timestamp 1713227210
<< nmos >>
rect -358 -81 -158 19
rect -100 -81 100 19
rect 158 -81 358 19
<< ndiff >>
rect -416 7 -358 19
rect -416 -69 -404 7
rect -370 -69 -358 7
rect -416 -81 -358 -69
rect -158 7 -100 19
rect -158 -69 -146 7
rect -112 -69 -100 7
rect -158 -81 -100 -69
rect 100 7 158 19
rect 100 -69 112 7
rect 146 -69 158 7
rect 100 -81 158 -69
rect 358 7 416 19
rect 358 -69 370 7
rect 404 -69 416 7
rect 358 -81 416 -69
<< ndiffc >>
rect -404 -69 -370 7
rect -146 -69 -112 7
rect 112 -69 146 7
rect 370 -69 404 7
<< poly >>
rect -358 91 -158 107
rect -358 57 -342 91
rect -174 57 -158 91
rect -358 19 -158 57
rect -100 91 100 107
rect -100 57 -84 91
rect 84 57 100 91
rect -100 19 100 57
rect 158 91 358 107
rect 158 57 174 91
rect 342 57 358 91
rect 158 19 358 57
rect -358 -107 -158 -81
rect -100 -107 100 -81
rect 158 -107 358 -81
<< polycont >>
rect -342 57 -174 91
rect -84 57 84 91
rect 174 57 342 91
<< locali >>
rect -358 57 -342 91
rect -174 57 -158 91
rect -100 57 -84 91
rect 84 57 100 91
rect 158 57 174 91
rect 342 57 358 91
rect -404 7 -370 23
rect -404 -85 -370 -69
rect -146 7 -112 23
rect -146 -85 -112 -69
rect 112 7 146 23
rect 112 -85 146 -69
rect 370 7 404 23
rect 370 -85 404 -69
<< viali >>
rect -342 57 -174 91
rect -84 57 84 91
rect 174 57 342 91
rect -404 -69 -370 7
rect -146 -69 -112 7
rect 112 -69 146 7
rect 370 -69 404 7
<< metal1 >>
rect -354 91 -162 97
rect -354 57 -342 91
rect -174 57 -162 91
rect -354 51 -162 57
rect -96 91 96 97
rect -96 57 -84 91
rect 84 57 96 91
rect -96 51 96 57
rect 162 91 354 97
rect 162 57 174 91
rect 342 57 354 91
rect 162 51 354 57
rect -410 7 -364 19
rect -410 -69 -404 7
rect -370 -69 -364 7
rect -410 -81 -364 -69
rect -152 7 -106 19
rect -152 -69 -146 7
rect -112 -69 -106 7
rect -152 -81 -106 -69
rect 106 7 152 19
rect 106 -69 112 7
rect 146 -69 152 7
rect 106 -81 152 -69
rect 364 7 410 19
rect 364 -69 370 7
rect 404 -69 410 7
rect 364 -81 410 -69
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.5 l 1 m 1 nf 3 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
