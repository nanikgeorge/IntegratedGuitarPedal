* NGSPICE file created from myOpamp.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_PE7Z8M a_1003_n64# a_1061_n161# a_n803_n64# a_n1319_n64#
+ a_1261_n64# a_n487_n161# a_n1261_n161# a_545_n161# a_745_n64# a_229_n64# w_n1355_n164#
+ a_n1061_n64# a_n545_n64# a_29_n161# a_487_n64# a_n745_n161# a_n29_n64# a_803_n161#
+ a_n287_n64# a_n229_n161# a_287_n161# a_n1003_n161# VSUBS
X0 a_n803_n64# a_n1003_n161# a_n1061_n64# w_n1355_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1 a_n29_n64# a_n229_n161# a_n287_n64# w_n1355_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2 a_745_n64# a_545_n161# a_487_n64# w_n1355_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3 a_229_n64# a_29_n161# a_n29_n64# w_n1355_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X4 a_487_n64# a_287_n161# a_229_n64# w_n1355_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X5 a_n545_n64# a_n745_n161# a_n803_n64# w_n1355_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X6 a_1261_n64# a_1061_n161# a_1003_n64# w_n1355_n164# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X7 a_n1061_n64# a_n1261_n161# a_n1319_n64# w_n1355_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X8 a_n287_n64# a_n487_n161# a_n545_n64# w_n1355_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X9 a_1003_n64# a_803_n161# a_745_n64# w_n1355_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
C0 w_n1355_n164# a_29_n161# 0.10872f
C1 a_545_n161# a_487_n64# 0.026809f
C2 a_287_n161# w_n1355_n164# 0.10872f
C3 a_745_n64# a_803_n161# 0.026809f
C4 a_n1061_n64# w_n1355_n164# 0.005183f
C5 w_n1355_n164# a_n229_n161# 0.10872f
C6 w_n1355_n164# a_n745_n161# 0.10872f
C7 w_n1355_n164# a_n1261_n161# 0.114821f
C8 a_745_n64# a_545_n161# 0.026809f
C9 a_n1061_n64# a_n1003_n161# 0.026809f
C10 a_n803_n64# a_n1061_n64# 0.055609f
C11 a_803_n161# a_545_n161# 0.061903f
C12 a_n1003_n161# a_n745_n161# 0.061903f
C13 a_n745_n161# a_n545_n64# 0.026809f
C14 a_n803_n64# a_n745_n161# 0.026809f
C15 a_n1003_n161# a_n1261_n161# 0.061903f
C16 a_487_n64# w_n1355_n164# 0.005183f
C17 a_n29_n64# a_29_n161# 0.026809f
C18 a_1061_n161# a_803_n161# 0.061903f
C19 w_n1355_n164# a_229_n64# 0.005183f
C20 a_287_n161# a_29_n161# 0.061903f
C21 a_n487_n161# a_n287_n64# 0.026809f
C22 a_n29_n64# a_n229_n161# 0.026809f
C23 a_745_n64# w_n1355_n164# 0.005183f
C24 a_n229_n161# a_29_n161# 0.061903f
C25 a_803_n161# w_n1355_n164# 0.10872f
C26 a_n1319_n64# w_n1355_n164# 0.008086f
C27 a_745_n64# a_1003_n64# 0.055609f
C28 w_n1355_n164# a_n487_n161# 0.10872f
C29 a_1003_n64# a_803_n161# 0.026809f
C30 a_545_n161# w_n1355_n164# 0.10872f
C31 a_n1061_n64# a_n1261_n161# 0.026809f
C32 a_487_n64# a_287_n161# 0.026809f
C33 a_n487_n161# a_n545_n64# 0.026809f
C34 w_n1355_n164# a_n287_n64# 0.005183f
C35 a_n29_n64# a_229_n64# 0.055609f
C36 a_1061_n161# w_n1355_n164# 0.114821f
C37 a_229_n64# a_29_n161# 0.026809f
C38 a_287_n161# a_229_n64# 0.026809f
C39 a_1061_n161# a_1261_n64# 0.026809f
C40 a_n545_n64# a_n287_n64# 0.055609f
C41 a_1061_n161# a_1003_n64# 0.026809f
C42 a_1261_n64# w_n1355_n164# 0.008086f
C43 a_n1319_n64# a_n1061_n64# 0.055609f
C44 w_n1355_n164# a_n1003_n161# 0.10872f
C45 a_1003_n64# w_n1355_n164# 0.005183f
C46 w_n1355_n164# a_n545_n64# 0.005183f
C47 a_n803_n64# w_n1355_n164# 0.005183f
C48 a_545_n161# a_287_n161# 0.061903f
C49 a_n29_n64# a_n287_n64# 0.055609f
C50 a_n487_n161# a_n229_n161# 0.061903f
C51 a_487_n64# a_229_n64# 0.055609f
C52 a_1003_n64# a_1261_n64# 0.055609f
C53 a_n1319_n64# a_n1261_n161# 0.026809f
C54 a_n487_n161# a_n745_n161# 0.061903f
C55 a_n803_n64# a_n1003_n161# 0.026809f
C56 a_745_n64# a_487_n64# 0.055609f
C57 a_n803_n64# a_n545_n64# 0.055609f
C58 a_n229_n161# a_n287_n64# 0.026809f
C59 a_n29_n64# w_n1355_n164# 0.005183f
C60 a_1261_n64# VSUBS 0.119027f
C61 a_1003_n64# VSUBS 0.051659f
C62 a_745_n64# VSUBS 0.051659f
C63 a_487_n64# VSUBS 0.051659f
C64 a_229_n64# VSUBS 0.051659f
C65 a_n29_n64# VSUBS 0.051659f
C66 a_n287_n64# VSUBS 0.051659f
C67 a_n545_n64# VSUBS 0.051659f
C68 a_n803_n64# VSUBS 0.051659f
C69 a_n1061_n64# VSUBS 0.051659f
C70 a_n1319_n64# VSUBS 0.119027f
C71 a_1061_n161# VSUBS 0.375556f
C72 a_803_n161# VSUBS 0.345228f
C73 a_545_n161# VSUBS 0.345228f
C74 a_287_n161# VSUBS 0.345228f
C75 a_29_n161# VSUBS 0.345228f
C76 a_n229_n161# VSUBS 0.345228f
C77 a_n487_n161# VSUBS 0.345228f
C78 a_n745_n161# VSUBS 0.345228f
C79 a_n1003_n161# VSUBS 0.345228f
C80 a_n1261_n161# VSUBS 0.375556f
C81 w_n1355_n164# VSUBS 2.94306f
.ends

.subckt sky130_fd_pr__nfet_01v8_7AMGGK a_n100_n157# a_n158_n69# a_100_n69# VSUBS
X0 a_100_n69# a_n100_n157# a_n158_n69# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
C0 a_n100_n157# a_100_n69# 0.026809f
C1 a_n100_n157# a_n158_n69# 0.026809f
C2 a_100_n69# a_n158_n69# 0.055609f
C3 a_100_n69# VSUBS 0.127112f
C4 a_n158_n69# VSUBS 0.127112f
C5 a_n100_n157# VSUBS 0.51752f
.ends

.subckt sky130_fd_pr__pfet_01v8_M2ZTWU a_n158_n64# w_n194_n164# a_n100_n161# a_100_n64#
+ VSUBS
X0 a_100_n64# a_n100_n161# a_n158_n64# w_n194_n164# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
C0 w_n194_n164# a_n158_n64# 0.008086f
C1 w_n194_n164# a_n100_n161# 0.120922f
C2 a_100_n64# w_n194_n164# 0.008086f
C3 a_n158_n64# a_n100_n161# 0.026809f
C4 a_100_n64# a_n158_n64# 0.055609f
C5 a_100_n64# a_n100_n161# 0.026809f
C6 a_100_n64# VSUBS 0.119027f
C7 a_n158_n64# VSUBS 0.119027f
C8 a_n100_n161# VSUBS 0.405884f
C9 w_n194_n164# VSUBS 0.421368f
.ends

.subckt sky130_fd_pr__nfet_01v8_HZNKM2 a_n229_n99# a_n545_n73# a_487_n73# a_n29_n73#
+ a_n487_n99# a_n287_n73# a_545_n99# a_29_n99# a_n803_n73# a_287_n99# a_745_n73# a_229_n73#
+ a_n745_n99# VSUBS
X0 a_n545_n73# a_n745_n99# a_n803_n73# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=1
X1 a_n287_n73# a_n487_n99# a_n545_n73# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X2 a_n29_n73# a_n229_n99# a_n287_n73# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X3 a_745_n73# a_545_n99# a_487_n73# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=1
X4 a_229_n73# a_29_n99# a_n29_n73# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X5 a_487_n73# a_287_n99# a_229_n73# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
C0 a_n229_n99# a_n29_n73# 0.014414f
C1 a_545_n99# a_487_n73# 0.014414f
C2 a_n803_n73# a_n545_n73# 0.02396f
C3 a_287_n99# a_487_n73# 0.014414f
C4 a_29_n99# a_n29_n73# 0.014414f
C5 a_29_n99# a_229_n73# 0.014414f
C6 a_n229_n99# a_n287_n73# 0.014414f
C7 a_n545_n73# a_n487_n99# 0.014414f
C8 a_n745_n99# a_n803_n73# 0.014414f
C9 a_229_n73# a_n29_n73# 0.02396f
C10 a_n287_n73# a_n487_n99# 0.014414f
C11 a_29_n99# a_287_n99# 0.05942f
C12 a_545_n99# a_745_n73# 0.014414f
C13 a_n29_n73# a_n287_n73# 0.02396f
C14 a_n745_n99# a_n487_n99# 0.05942f
C15 a_229_n73# a_287_n99# 0.014414f
C16 a_745_n73# a_487_n73# 0.02396f
C17 a_n545_n73# a_n287_n73# 0.02396f
C18 a_n229_n99# a_n487_n99# 0.05942f
C19 a_287_n99# a_545_n99# 0.05942f
C20 a_29_n99# a_n229_n99# 0.05942f
C21 a_229_n73# a_487_n73# 0.02396f
C22 a_n745_n99# a_n545_n73# 0.014414f
C23 a_745_n73# VSUBS 0.072287f
C24 a_487_n73# VSUBS 0.041002f
C25 a_229_n73# VSUBS 0.041002f
C26 a_n29_n73# VSUBS 0.041002f
C27 a_n287_n73# VSUBS 0.041002f
C28 a_n545_n73# VSUBS 0.041002f
C29 a_n803_n73# VSUBS 0.072287f
C30 a_545_n99# VSUBS 0.489687f
C31 a_287_n99# VSUBS 0.454871f
C32 a_29_n99# VSUBS 0.454871f
C33 a_n229_n99# VSUBS 0.454871f
C34 a_n487_n99# VSUBS 0.454871f
C35 a_n745_n99# VSUBS 0.489687f
.ends

.subckt sky130_fd_pr__nfet_01v8_DVNKMG a_158_n99# a_100_n73# a_n100_n99# a_n416_n73#
+ a_358_n73# a_n358_n99# a_n158_n73# VSUBS
X0 a_358_n73# a_158_n99# a_100_n73# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=1
X1 a_n158_n73# a_n358_n99# a_n416_n73# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=1
X2 a_100_n73# a_n100_n99# a_n158_n73# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
C0 a_358_n73# a_158_n99# 0.014414f
C1 a_n358_n99# a_n100_n99# 0.05942f
C2 a_n158_n73# a_n416_n73# 0.02396f
C3 a_n158_n73# a_100_n73# 0.02396f
C4 a_n100_n99# a_100_n73# 0.014414f
C5 a_158_n99# a_100_n73# 0.014414f
C6 a_n158_n73# a_n100_n99# 0.014414f
C7 a_358_n73# a_100_n73# 0.02396f
C8 a_n100_n99# a_158_n99# 0.05942f
C9 a_n358_n99# a_n416_n73# 0.014414f
C10 a_n158_n73# a_n358_n99# 0.014414f
C11 a_358_n73# VSUBS 0.072287f
C12 a_100_n73# VSUBS 0.041002f
C13 a_n158_n73# VSUBS 0.041002f
C14 a_n416_n73# VSUBS 0.072287f
C15 a_158_n99# VSUBS 0.489687f
C16 a_n100_n99# VSUBS 0.454871f
C17 a_n358_n99# VSUBS 0.489687f
.ends

.subckt sky130_fd_pr__nfet_01v8_QFRGQ5 a_100_n131# a_n100_n157# a_n158_n131# VSUBS
X0 a_100_n131# a_n100_n157# a_n158_n131# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
C0 a_100_n131# a_n158_n131# 0.055609f
C1 a_n158_n131# a_n100_n157# 0.026809f
C2 a_100_n131# a_n100_n157# 0.026809f
C3 a_100_n131# VSUBS 0.127112f
C4 a_n158_n131# VSUBS 0.127112f
C5 a_n100_n157# VSUBS 0.51752f
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_JNUKDP a_546_n568# a_n616_n568# VSUBS
X0 a_546_n568# a_n616_n568# VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=26.11
C0 a_546_n568# a_n616_n568# 0.019671f
C1 a_546_n568# VSUBS 0.395178f
C2 a_n616_n568# VSUBS 0.395178f
.ends

.subckt sky130_fd_pr__nfet_01v8_2F8GYT a_n100_n157# a_n158_n69# a_100_n69# VSUBS
X0 a_100_n69# a_n100_n157# a_n158_n69# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
C0 a_100_n69# a_n158_n69# 0.055609f
C1 a_n158_n69# a_n100_n157# 0.026809f
C2 a_100_n69# a_n100_n157# 0.026809f
C3 a_100_n69# VSUBS 0.127112f
C4 a_n158_n69# VSUBS 0.127112f
C5 a_n100_n157# VSUBS 0.51752f
.ends

.subckt myOpamp VDD OUT INp INn VSS
Xsky130_fd_pr__pfet_01v8_PE7Z8M_0 VDD m1_280_190# OUT m1_280_190# OUT m1_280_190#
+ m1_280_190# m1_280_190# m1_280_190# OUT VDD VDD VDD m1_280_190# VDD m1_280_190#
+ VDD m1_280_190# m1_280_190# m1_280_190# m1_280_190# m1_280_190# VSS sky130_fd_pr__pfet_01v8_PE7Z8M
Xsky130_fd_pr__nfet_01v8_7AMGGK_0 INn m1_540_190# OUT VSS sky130_fd_pr__nfet_01v8_7AMGGK
Xsky130_fd_pr__nfet_01v8_7AMGGK_1 INn OUT m1_540_190# VSS sky130_fd_pr__nfet_01v8_7AMGGK
Xsky130_fd_pr__nfet_01v8_7AMGGK_3 INn m1_540_190# OUT VSS sky130_fd_pr__nfet_01v8_7AMGGK
Xsky130_fd_pr__nfet_01v8_7AMGGK_4 INn m1_540_190# OUT VSS sky130_fd_pr__nfet_01v8_7AMGGK
Xsky130_fd_pr__nfet_01v8_7AMGGK_5 INn OUT m1_540_190# VSS sky130_fd_pr__nfet_01v8_7AMGGK
Xsky130_fd_pr__pfet_01v8_M2ZTWU_0 VDD VDD VDD m1_280_190# VSS sky130_fd_pr__pfet_01v8_M2ZTWU
Xsky130_fd_pr__nfet_01v8_HZNKM2_0 li_n480_n300# m1_540_190# m1_540_190# li_n480_n300#
+ li_n480_n300# VSS li_n480_n300# li_n480_n300# VSS li_n480_n300# VSS VSS li_n480_n300#
+ VSS sky130_fd_pr__nfet_01v8_HZNKM2
Xsky130_fd_pr__nfet_01v8_DVNKMG_0 VSS VSS VSS VSS VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_DVNKMG
Xsky130_fd_pr__pfet_01v8_M2ZTWU_1 OUT VDD VDD VDD VSS sky130_fd_pr__pfet_01v8_M2ZTWU
Xsky130_fd_pr__nfet_01v8_DVNKMG_1 VSS VSS VSS VSS VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_DVNKMG
Xsky130_fd_pr__nfet_01v8_QFRGQ5_0 m1_540_190# INp m1_280_190# VSS sky130_fd_pr__nfet_01v8_QFRGQ5
Xsky130_fd_pr__nfet_01v8_QFRGQ5_1 m1_280_190# INp m1_540_190# VSS sky130_fd_pr__nfet_01v8_QFRGQ5
Xsky130_fd_pr__nfet_01v8_QFRGQ5_2 m1_540_190# INp m1_280_190# VSS sky130_fd_pr__nfet_01v8_QFRGQ5
Xsky130_fd_pr__res_xhigh_po_0p35_JNUKDP_0 VDD li_n480_n300# VSS sky130_fd_pr__res_xhigh_po_0p35_JNUKDP
Xsky130_fd_pr__nfet_01v8_QFRGQ5_3 m1_280_190# INp m1_540_190# VSS sky130_fd_pr__nfet_01v8_QFRGQ5
Xsky130_fd_pr__nfet_01v8_QFRGQ5_5 m1_540_190# INp m1_280_190# VSS sky130_fd_pr__nfet_01v8_QFRGQ5
Xsky130_fd_pr__nfet_01v8_2F8GYT_0 VSS OUT VSS VSS sky130_fd_pr__nfet_01v8_2F8GYT
Xsky130_fd_pr__nfet_01v8_2F8GYT_1 VSS VSS m1_280_190# VSS sky130_fd_pr__nfet_01v8_2F8GYT
C0 VDD VSS 0.132689f
C1 li_n480_n300# VSS 0.543414f
C2 m1_280_190# OUT 2.216533f
C3 INn OUT 0.897128f
C4 m1_540_190# VDD 0.137313f
C5 INn m1_280_190# 0.8459f
C6 m1_540_190# li_n480_n300# 1.474142f
C7 INp VDD 0.673697f
C8 li_n480_n300# INp 0.162656f
C9 m1_540_190# VSS -0.030498f
C10 INp VSS 0.12778f
C11 OUT VDD 1.608392f
C12 li_n480_n300# OUT 0.001336f
C13 m1_280_190# VDD 2.650126f
C14 INn VDD 0.172036f
C15 li_n480_n300# m1_280_190# 0.275219f
C16 li_n480_n300# INn 1.130703f
C17 m1_540_190# INp 0.626583f
C18 OUT VSS -0.017714f
C19 m1_280_190# VSS 0.015251f
C20 INn VSS 0.277875f
C21 m1_540_190# OUT 0.383989f
C22 li_n480_n300# VDD 0.077209f
C23 m1_540_190# m1_280_190# 1.299842f
C24 m1_540_190# INn 1.100506f
C25 INp OUT 0.763432f
C26 m1_280_190# INp 2.951741f
C27 INn INp 0.499442f
C28 m1_540_190# 0 1.525095f
C29 m1_280_190# 0 2.597431f
C30 INp 0 1.663726f
C31 VSS 0 1.6306f
C32 li_n480_n300# 0 4.729789f
C33 OUT 0 0.416294f
C34 INn 0 2.23613f
C35 VDD 0 40.724533f
.ends

