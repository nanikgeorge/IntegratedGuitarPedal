magic
tech sky130A
magscale 1 2
timestamp 1712972901
<< error_p >>
rect -31 145 31 151
rect -31 111 -19 145
rect -31 105 31 111
<< nwell >>
rect -129 -198 129 164
<< pmos >>
rect -35 -136 35 64
<< pdiff >>
rect -93 52 -35 64
rect -93 -124 -81 52
rect -47 -124 -35 52
rect -93 -136 -35 -124
rect 35 52 93 64
rect 35 -124 47 52
rect 81 -124 93 52
rect 35 -136 93 -124
<< pdiffc >>
rect -81 -124 -47 52
rect 47 -124 81 52
<< poly >>
rect -35 145 35 161
rect -35 111 -19 145
rect 19 111 35 145
rect -35 64 35 111
rect -35 -162 35 -136
<< polycont >>
rect -19 111 19 145
<< locali >>
rect -35 111 -19 145
rect 19 111 35 145
rect -81 52 -47 68
rect -81 -140 -47 -124
rect 47 52 81 68
rect 47 -140 81 -124
<< viali >>
rect -19 111 19 145
rect -81 -124 -47 52
rect 47 -124 81 52
<< metal1 >>
rect -31 145 31 151
rect -31 111 -19 145
rect 19 111 31 145
rect -31 105 31 111
rect -87 52 -41 64
rect -87 -124 -81 52
rect -47 -124 -41 52
rect -87 -136 -41 -124
rect 41 52 87 64
rect 41 -124 47 52
rect 81 -124 87 52
rect 41 -136 87 -124
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.35 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
