* NGSPICE file created from distortion_flat2.ext - technology: sky130A
*IN VSS OUT CTRL VDD
.subckt distortion_unit VDD CTRL IN OUT VSS
X0 a_1740_1605# a_1740_1605# VDD.t35 VDD.t34 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1 VDD.t33 a_1740_1605# tgate_1.IN VDD.t32 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2 tgate_1.IN a_1740_1605# VDD.t31 VDD.t30 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3 a_1740_1605# IN.t4 a_1998_1605# VSS.t46 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X4 a_1998_1605# IN.t5 a_1740_1605# VSS.t45 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X5 tgate_0.CTRL CTRL.t0 VDD.t38 sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VSS.t55 a_944_1150# a_1998_1605# VSS.t44 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X7 VDD.t9 CTRL.t1 tgate_0.CTRL sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8 a_1998_1605# a_944_1150# VSS.t54 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X9 VDD.t36 CTRL.t2 tgate_0.CTRL sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VSS.t53 a_944_1150# a_944_1150# VSS.t37 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X11 tgate_0.CTRL CTRL.t3 VDD.t2 sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 VDD.t8 a_944_1150# VSS.t43 sky130_fd_pr__res_xhigh_po_0p35 l=0.16
X13 tgate_0.CTRL CTRL.t4 VDD.t1 sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X14 tgate_0.CTRL CTRL.t5 VSS.t6 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VDD.t29 a_1740_1605# a_1740_1605# VDD.t28 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X16 tgate_1.IN tgate_0.CTRL OUT.t5 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X17 a_1740_1605# VDD.t13 VDD.t15 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X18 VDD.t27 a_1740_1605# a_1740_1605# VDD.t26 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X19 VDD.t37 CTRL.t6 tgate_0.CTRL sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 a_1740_1605# IN.t6 a_1998_1605# VSS.t44 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X21 VSS.t35 VSS.t33 VSS.t35 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X22 OUT.t1 CTRL.t7 tgate_1.IN VSS.t57 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X23 VSS.t4 CTRL.t8 tgate_0.CTRL VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 OUT.t3 CTRL.t9 IN.t3 VDD.t7 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X25 a_1998_1605# myOpamp_0.INn tgate_1.IN VSS.t38 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X26 VSS.t32 VSS.t30 VSS.t31 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0 ps=0 w=0.42 l=1
X27 VSS.t29 VSS.t27 VSS.t29 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X28 tgate_1.IN myOpamp_0.INn a_1998_1605# VSS.t37 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X29 IN.t1 tgate_0.CTRL OUT.t7 VSS.t40 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X30 a_3626_n94# myOpamp_0.INn VSS.t49 sky130_fd_pr__res_xhigh_po_0p35 l=4
X31 tgate_1.IN myOpamp_0.INn VSS.t56 sky130_fd_pr__res_xhigh_po_0p35 l=10
X32 tgate_0.CTRL CTRL.t10 VSS.t2 VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X33 VDD.t25 a_1740_1605# tgate_1.IN VDD.t24 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X34 VDD.t12 VDD.t10 tgate_1.IN VDD.t11 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X35 tgate_0.CTRL CTRL.t11 VSS.t10 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X36 tgate_1.IN a_1740_1605# VDD.t23 VDD.t22 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X37 tgate_1.IN a_1740_1605# VDD.t21 VDD.t20 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X38 a_1740_1605# VSS.t24 VSS.t26 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X39 a_1998_1605# IN.t7 a_1740_1605# VSS.t34 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X40 a_1998_1605# IN.t8 a_1740_1605# VSS.t28 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X41 a_1998_1605# a_944_1150# VSS.t52 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X42 VSS.t23 VSS.t22 VSS.t23 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X43 tgate_0.CTRL CTRL.t12 VDD.t3 sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X44 VSS.t21 VSS.t19 VSS.t21 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X45 VSS.t18 VSS.t16 VSS.t18 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X46 OUT.t4 tgate_0.CTRL tgate_1.IN VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X47 tgate_0.CTRL CTRL.t13 VSS.t12 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X48 a_1740_1605# a_1740_1605# VDD.t19 VDD.t18 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X49 VDD.t17 a_1740_1605# a_1740_1605# VDD.t16 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X50 tgate_1.IN CTRL.t14 OUT.t0 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X51 VSS.t48 CTRL.t15 tgate_0.CTRL VSS.t47 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X52 a_1998_1605# myOpamp_0.INn tgate_1.IN VSS.t36 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X53 VSS.t15 VSS.t13 tgate_1.IN VSS.t14 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X54 VSS.t51 a_944_1150# a_1998_1605# VSS.t46 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X55 a_944_1150# a_944_1150# VSS.t50 VSS.t45 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X56 tgate_1.IN myOpamp_0.INn a_1998_1605# VSS.t20 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X57 tgate_1.IN myOpamp_0.INn a_1998_1605# VSS.t17 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X58 IN.t0 CTRL.t16 OUT.t2 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X59 VDD a_944_1150# VSS sky130_fd_pr__res_xhigh_po_0p35 l=26.11
X60 VDD.t4 CTRL.t17 tgate_0.CTRL sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X61 VSS.t42 CTRL.t18 tgate_0.CTRL VSS.t41 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X62 OUT.t6 tgate_0.CTRL IN.t2 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X63 VSS.t8 CTRL.t19 tgate_0.CTRL VSS.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 VDD.n14 VDD.n13 18810
R1 VDD.n15 VDD.n14 18786.2
R2 VDD.n15 VDD.n6 18786.2
R3 VDD.n13 VDD.n6 18667.5
R4 VDD.n16 VDD.n4 7334.54
R5 VDD.n12 VDD.n5 7332.73
R6 VDD.n16 VDD.n5 7312.73
R7 VDD.n12 VDD.n4 7300
R8 VDD.n41 VDD.n39 4136.47
R9 VDD.n48 VDD.n46 4136.47
R10 VDD.n41 VDD.n38 2068.24
R11 VDD.n48 VDD.n45 2068.24
R12 VDD.n10 VDD.n8 781.188
R13 VDD.n18 VDD.n2 779.442
R14 VDD.n17 VDD.n3 779.056
R15 VDD.n11 VDD.n7 778.668
R16 VDD.t20 VDD.t11 478.712
R17 VDD.t26 VDD.t20 478.712
R18 VDD.t34 VDD.t26 478.712
R19 VDD.t32 VDD.t34 478.712
R20 VDD.t30 VDD.t32 478.712
R21 VDD.t16 VDD.t18 478.712
R22 VDD.t18 VDD.t24 478.712
R23 VDD.t24 VDD.t22 478.712
R24 VDD.t22 VDD.t28 478.712
R25 VDD.t28 VDD.t14 478.712
R26 VDD.n41 VDD.t0 452.676
R27 VDD.t7 VDD.n39 452.676
R28 VDD.n48 VDD.t6 452.676
R29 VDD.t5 VDD.n46 452.676
R30 VDD.n67 VDD.t1 342.377
R31 VDD.n57 VDD.t9 338.892
R32 VDD.n72 VDD.n65 320.976
R33 VDD.n64 VDD.n54 320.976
R34 VDD.n62 VDD.n55 320.976
R35 VDD.n31 VDD.t16 269.043
R36 VDD.n32 VDD.t8 264.031
R37 VDD.n26 VDD.t15 228.215
R38 VDD.n21 VDD.t12 228.215
R39 VDD.t0 VDD.n40 215.757
R40 VDD.n40 VDD.t7 215.757
R41 VDD.t6 VDD.n47 215.757
R42 VDD.n47 VDD.t5 215.757
R43 VDD.n31 VDD.t30 209.668
R44 VDD.n28 VDD.n27 199.851
R45 VDD.n30 VDD.n29 199.851
R46 VDD.n23 VDD.n22 199.851
R47 VDD.n25 VDD.n24 199.851
R48 VDD.n35 VDD.n34 199.851
R49 VDD.n39 VDD.n37 163.684
R50 VDD.n46 VDD.n44 163.684
R51 VDD.n21 VDD.t10 120.855
R52 VDD.n26 VDD.t13 120.749
R53 VDD.n42 VDD.n37 113.915
R54 VDD.n49 VDD.n44 113.915
R55 VDD.n42 VDD.n41 47.0382
R56 VDD.n49 VDD.n48 47.0382
R57 VDD.n32 VDD.n31 38.8096
R58 VDD.n57 VDD 35.5709
R59 VDD.n61 VDD.n56 34.6358
R60 VDD.n74 VDD.n73 34.6358
R61 VDD.n71 VDD.n66 34.6358
R62 VDD.n64 VDD.n63 32.0005
R63 VDD.n63 VDD.n62 31.2476
R64 VDD.n27 VDD.t23 28.5655
R65 VDD.n27 VDD.t29 28.5655
R66 VDD.n29 VDD.t19 28.5655
R67 VDD.n29 VDD.t25 28.5655
R68 VDD.n22 VDD.t21 28.5655
R69 VDD.n22 VDD.t27 28.5655
R70 VDD.n24 VDD.t35 28.5655
R71 VDD.n24 VDD.t33 28.5655
R72 VDD.n34 VDD.t31 28.5655
R73 VDD.n34 VDD.t17 28.5655
R74 VDD.n65 VDD.t38 26.5955
R75 VDD.n65 VDD.t36 26.5955
R76 VDD.n54 VDD.t3 26.5955
R77 VDD.n54 VDD.t4 26.5955
R78 VDD.n55 VDD.t2 26.5955
R79 VDD.n55 VDD.t37 26.5955
R80 VDD.n73 VDD.n72 25.977
R81 VDD.n40 VDD.n38 20.5561
R82 VDD.n47 VDD.n45 20.5561
R83 VDD.n57 VDD.n56 18.824
R84 VDD.n38 VDD.n37 18.7435
R85 VDD.n45 VDD.n44 18.7435
R86 VDD.n67 VDD.n66 13.5534
R87 VDD VDD.n42 11.4981
R88 VDD VDD.n49 11.4981
R89 VDD.n68 VDD.n67 11.1829
R90 VDD.n58 VDD.n57 9.3005
R91 VDD.n59 VDD.n56 9.3005
R92 VDD.n61 VDD.n60 9.3005
R93 VDD.n63 VDD.n52 9.3005
R94 VDD.n75 VDD.n74 9.3005
R95 VDD.n73 VDD.n53 9.3005
R96 VDD.n71 VDD.n70 9.3005
R97 VDD.n69 VDD.n66 9.3005
R98 VDD.n72 VDD.n71 8.65932
R99 VDD.n8 VDD.n5 5.0005
R100 VDD.n14 VDD.n5 5.0005
R101 VDD.n7 VDD.n4 4.86892
R102 VDD.n6 VDD.n4 4.86892
R103 VDD.n62 VDD.n61 3.38874
R104 VDD.n51 VDD.n50 3.28283
R105 VDD.n51 VDD.n43 3.19667
R106 VDD.n74 VDD.n64 2.63579
R107 VDD.n19 VDD.n1 2.4755
R108 VDD.n9 VDD.n1 2.4755
R109 VDD.n9 VDD.n0 2.463
R110 VDD.n17 VDD.n16 2.34227
R111 VDD.n16 VDD.n15 2.34227
R112 VDD.n12 VDD.n11 2.34227
R113 VDD.n13 VDD.n12 2.34227
R114 VDD.n20 VDD.n0 2.10363
R115 VDD.n18 VDD.n17 1.93989
R116 VDD.n77 VDD.n76 1.02714
R117 VDD.n7 VDD.n2 0.970197
R118 VDD.n11 VDD.n10 0.970197
R119 VDD.n8 VDD.n3 0.970197
R120 VDD.n23 VDD.n21 0.890989
R121 VDD.n28 VDD.n26 0.760446
R122 VDD.n77 VDD.n51 0.419651
R123 VDD.n30 VDD.n28 0.40675
R124 VDD.n25 VDD.n23 0.40675
R125 VDD.n35 VDD.n25 0.40675
R126 VDD.n20 VDD.n19 0.359875
R127 VDD.n3 VDD.n1 0.258833
R128 VDD.n2 VDD.n0 0.258833
R129 VDD.n78 VDD.n77 0.257907
R130 VDD.n35 VDD.n33 0.208833
R131 VDD.n33 VDD.n30 0.188
R132 VDD.n33 VDD.n32 0.1865
R133 VDD.n78 VDD 0.15243
R134 VDD.n10 VDD.n9 0.121279
R135 VDD.n19 VDD.n18 0.121279
R136 VDD.n59 VDD.n58 0.120292
R137 VDD.n60 VDD.n59 0.120292
R138 VDD.n60 VDD.n52 0.120292
R139 VDD.n75 VDD.n53 0.120292
R140 VDD.n70 VDD.n53 0.120292
R141 VDD.n70 VDD.n69 0.120292
R142 VDD.n69 VDD.n68 0.120292
R143 VDD.n76 VDD.n75 0.115083
R144 VDD VDD.n80 0.096686
R145 VDD.n36 VDD.n35 0.0948367
R146 VDD.n36 VDD.n20 0.0691538
R147 VDD.n79 VDD.n36 0.0614341
R148 VDD.n58 VDD 0.0603958
R149 VDD VDD.n79 0.0562442
R150 VDD.n43 VDD 0.0459545
R151 VDD.n50 VDD 0.0459545
R152 VDD.n43 VDD 0.0338333
R153 VDD.n50 VDD 0.0338333
R154 VDD.n68 VDD 0.0226354
R155 VDD.n79 VDD.n78 0.00599114
R156 VDD.n76 VDD.n52 0.00570833
R157 IN.n4 IN.t0 223.565
R158 IN.n7 IN.t3 223.565
R159 IN.n0 IN.t8 118.769
R160 IN.n3 IN.t7 118.621
R161 IN.n2 IN.t4 118.005
R162 IN.n1 IN.t5 118.005
R163 IN.n0 IN.t6 118.005
R164 IN.n6 IN.n5 90.2112
R165 IN.n6 IN.n4 66.2405
R166 IN.n7 IN.n6 63.2157
R167 IN.n5 IN.t2 17.4005
R168 IN.n5 IN.t1 17.4005
R169 IN.n8 IN.n4 5.54823
R170 IN.n8 IN.n7 5.18686
R171 IN.n9 IN 4.4438
R172 IN IN.n3 2.77717
R173 IN.n1 IN.n0 2.66195
R174 IN.n3 IN.n2 1.71868
R175 IN.n2 IN.n1 0.764886
R176 IN IN.n9 0.490406
R177 IN IN.n8 0.244818
R178 IN.n9 IN 0.0129412
R179 VSS.n84 VSS.n83 80833
R180 VSS.n61 VSS.n60 27500
R181 VSS.n61 VSS.t43 10325.8
R182 VSS.n73 VSS.n55 10285.8
R183 VSS.n62 VSS.n55 10253
R184 VSS.n73 VSS.n56 10250
R185 VSS.n62 VSS.n56 10187.3
R186 VSS.n25 VSS.n23 9618.24
R187 VSS.n82 VSS.n23 9618.24
R188 VSS.n25 VSS.n17 9618.24
R189 VSS.n82 VSS.n17 9618.24
R190 VSS.n96 VSS.n6 9562.45
R191 VSS.n84 VSS.t49 7047.59
R192 VSS.n100 VSS.n3 6732.76
R193 VSS.n94 VSS.t49 6660.69
R194 VSS.n92 VSS.n5 6309.89
R195 VSS.n90 VSS.n18 6141.76
R196 VSS.n85 VSS.n18 6141.76
R197 VSS.n90 VSS.n19 6141.76
R198 VSS.n85 VSS.n19 6141.76
R199 VSS.n6 VSS.n5 4126.19
R200 VSS.n100 VSS.n4 3366.38
R201 VSS.n95 VSS.n94 2126.67
R202 VSS.n9 VSS.n7 1683.19
R203 VSS.n14 VSS.n7 1683.19
R204 VSS.t47 VSS.n92 1511.05
R205 VSS.n60 VSS.t14 1302.55
R206 VSS.t39 VSS.n10 1198.65
R207 VSS.n15 VSS.t40 1198.65
R208 VSS.n99 VSS.t57 1053.4
R209 VSS.t0 VSS.n97 1053.4
R210 VSS.n96 VSS.n95 967.52
R211 VSS.n12 VSS.n7 841.596
R212 VSS.n91 VSS.n17 835.168
R213 VSS.t14 VSS.t17 803.966
R214 VSS.t17 VSS.t28 803.966
R215 VSS.t28 VSS.t44 803.966
R216 VSS.t44 VSS.t38 803.966
R217 VSS.t38 VSS.t37 803.966
R218 VSS.t45 VSS.t46 803.966
R219 VSS.t20 VSS.t36 803.966
R220 VSS.t34 VSS.t20 803.966
R221 VSS.t25 VSS.t34 803.966
R222 VSS VSS.t11 785.428
R223 VSS.t9 VSS.t47 673.225
R224 VSS.t3 VSS.t9 673.225
R225 VSS.t1 VSS.t3 673.225
R226 VSS.t7 VSS.t1 673.225
R227 VSS.t5 VSS.t7 673.225
R228 VSS.t41 VSS.t5 673.225
R229 VSS.t11 VSS.t41 673.225
R230 VSS.n66 VSS.n57 666.376
R231 VSS.n72 VSS.n71 665.019
R232 VSS.n65 VSS.n64 664.242
R233 VSS.n63 VSS.n58 661.915
R234 VSS.t43 VSS.t25 660.674
R235 VSS.n11 VSS.t39 636.323
R236 VSS.n11 VSS.t40 636.323
R237 VSS.t46 VSS.n74 629.462
R238 VSS.n26 VSS.n24 624.942
R239 VSS.n27 VSS.n26 624.942
R240 VSS.n81 VSS.n27 624.942
R241 VSS.t57 VSS.n98 559.212
R242 VSS.n98 VSS.t0 559.212
R243 VSS.n93 VSS 536.976
R244 VSS.n92 VSS 469.406
R245 VSS.n75 VSS.t37 414.449
R246 VSS.n87 VSS.n86 399.757
R247 VSS.n88 VSS.n87 398.683
R248 VSS.n75 VSS.t45 389.519
R249 VSS.n89 VSS.n20 333.26
R250 VSS.n80 VSS.n21 314.127
R251 VSS.n86 VSS.n85 292.5
R252 VSS.n85 VSS.n84 292.5
R253 VSS.n27 VSS.n23 292.5
R254 VSS.n23 VSS.t56 292.5
R255 VSS.n90 VSS.n89 292.5
R256 VSS.n91 VSS.n90 292.5
R257 VSS.n24 VSS.n17 292.5
R258 VSS.n118 VSS.t12 287.151
R259 VSS.n107 VSS.t48 284.024
R260 VSS.n93 VSS.n91 267.668
R261 VSS.n10 VSS.n6 261.435
R262 VSS.n96 VSS.n15 261.435
R263 VSS.n14 VSS.n13 254.685
R264 VSS.n47 VSS.t32 236.113
R265 VSS.t23 VSS.n31 235.764
R266 VSS.n3 VSS.n2 232.597
R267 VSS.n99 VSS.n5 229.755
R268 VSS.n97 VSS.n96 229.755
R269 VSS.n112 VSS.n106 207.213
R270 VSS.n125 VSS.n113 207.213
R271 VSS.n115 VSS.n114 207.213
R272 VSS.n52 VSS.n51 194.805
R273 VSS.n38 VSS.n37 194.542
R274 VSS.n54 VSS.n53 194.463
R275 VSS.n40 VSS.n39 194.463
R276 VSS.n48 VSS.n47 194.3
R277 VSS.n50 VSS.n49 194.3
R278 VSS.n36 VSS.n35 194.3
R279 VSS.n33 VSS.n32 194.3
R280 VSS.n60 VSS.n55 189.166
R281 VSS.n83 VSS.t56 177.44
R282 VSS.n74 VSS.t36 174.505
R283 VSS.t56 VSS.n16 161.225
R284 VSS.n9 VSS.n8 147.038
R285 VSS.n101 VSS.n100 147.038
R286 VSS.n10 VSS.n9 146.25
R287 VSS.n15 VSS.n14 146.25
R288 VSS.n97 VSS.n3 146.25
R289 VSS.n100 VSS.n99 146.25
R290 VSS.n44 VSS.t24 118.005
R291 VSS.n30 VSS.t13 118.005
R292 VSS.n86 VSS.n22 111.401
R293 VSS.n24 VSS.n21 104.659
R294 VSS.n45 VSS.t30 104.028
R295 VSS.n43 VSS.t33 104.028
R296 VSS.n42 VSS.t19 104.028
R297 VSS.n28 VSS.t27 104.028
R298 VSS.n34 VSS.t16 104.028
R299 VSS.n29 VSS.t22 104.028
R300 VSS.n101 VSS.n2 92.9264
R301 VSS.n13 VSS.n8 88.4348
R302 VSS.n44 VSS.t26 87.6949
R303 VSS.n30 VSS.t15 87.5315
R304 VSS.n95 VSS.n16 77.3449
R305 VSS.t43 VSS.n56 77.0353
R306 VSS.n81 VSS.n80 66.4099
R307 VSS.n13 VSS.n12 65.0005
R308 VSS.n12 VSS.n11 65.0005
R309 VSS.n98 VSS.n4 65.0005
R310 VSS.n4 VSS.n2 59.3637
R311 VSS.n94 VSS.n93 58.6672
R312 VSS.n51 VSS.t52 41.4291
R313 VSS.n51 VSS.t21 41.4291
R314 VSS.t35 VSS.n48 41.4291
R315 VSS.n48 VSS.t31 41.4291
R316 VSS.t21 VSS.n50 41.4291
R317 VSS.n50 VSS.t35 41.4291
R318 VSS.n53 VSS.t50 41.4291
R319 VSS.n53 VSS.t51 41.4291
R320 VSS.n37 VSS.t29 41.4291
R321 VSS.n37 VSS.t55 41.4291
R322 VSS.n36 VSS.t18 41.4291
R323 VSS.t29 VSS.n36 41.4291
R324 VSS.n32 VSS.t23 41.4291
R325 VSS.n32 VSS.t18 41.4291
R326 VSS.n39 VSS.t54 41.4291
R327 VSS.n39 VSS.t53 41.4291
R328 VSS VSS.n107 35.197
R329 VSS.n111 VSS.n110 34.6358
R330 VSS.n124 VSS.n123 34.6358
R331 VSS.n120 VSS.n119 34.6358
R332 VSS.n22 VSS.n20 34.2005
R333 VSS.n126 VSS.n125 32.0005
R334 VSS.n126 VSS.n112 31.2476
R335 VSS.n76 VSS.n75 26.2219
R336 VSS.n123 VSS.n115 25.977
R337 VSS.n106 VSS.t10 24.9236
R338 VSS.n106 VSS.t4 24.9236
R339 VSS.n113 VSS.t2 24.9236
R340 VSS.n113 VSS.t8 24.9236
R341 VSS.n114 VSS.t6 24.9236
R342 VSS.n114 VSS.t42 24.9236
R343 VSS.n87 VSS.n19 23.4005
R344 VSS.n19 VSS.t49 23.4005
R345 VSS.n20 VSS.n18 23.4005
R346 VSS.n18 VSS.t49 23.4005
R347 VSS.n58 VSS.n56 20.8934
R348 VSS.n65 VSS.n55 20.8934
R349 VSS.n25 VSS.n16 18.8625
R350 VSS.n110 VSS.n107 18.824
R351 VSS.n82 VSS.n81 13.6052
R352 VSS.n83 VSS.n82 13.6052
R353 VSS.n26 VSS.n25 13.6052
R354 VSS.n119 VSS.n118 13.5534
R355 VSS.n8 VSS 11.4981
R356 VSS VSS.n101 11.4981
R357 VSS.n118 VSS.n117 11.1829
R358 VSS.n108 VSS.n107 9.3005
R359 VSS.n110 VSS.n109 9.3005
R360 VSS.n111 VSS.n104 9.3005
R361 VSS.n127 VSS.n126 9.3005
R362 VSS.n124 VSS.n105 9.3005
R363 VSS.n123 VSS.n122 9.3005
R364 VSS.n121 VSS.n120 9.3005
R365 VSS.n119 VSS.n116 9.3005
R366 VSS.n120 VSS.n115 8.65932
R367 VSS.n63 VSS.n62 8.23994
R368 VSS.n62 VSS.n61 8.23994
R369 VSS.n73 VSS.n72 8.23994
R370 VSS.n74 VSS.n73 8.23994
R371 VSS.n88 VSS.n21 5.9205
R372 VSS.n103 VSS.n1 3.45067
R373 VSS.n112 VSS.n111 3.38874
R374 VSS.n103 VSS.n102 2.87883
R375 VSS.n125 VSS.n124 2.63579
R376 VSS.n80 VSS.n79 2.45057
R377 VSS.n70 VSS.n59 2.09737
R378 VSS.n70 VSS.n69 2.09737
R379 VSS.n67 VSS.n59 2.09113
R380 VSS.n64 VSS.n63 1.93989
R381 VSS.n68 VSS.n67 1.72862
R382 VSS.n129 VSS.n128 1.24162
R383 VSS.n71 VSS.n58 0.970197
R384 VSS.n72 VSS.n57 0.970197
R385 VSS.n66 VSS.n65 0.970197
R386 VSS.n54 VSS.n52 0.927299
R387 VSS.n79 VSS.n22 0.846456
R388 VSS.n40 VSS.n38 0.690273
R389 VSS.n129 VSS.n103 0.6315
R390 VSS.n52 VSS.n41 0.60675
R391 VSS.n52 VSS.n46 0.516045
R392 VSS.n42 VSS.n41 0.454213
R393 VSS.n89 VSS.n88 0.376971
R394 VSS.n69 VSS.n68 0.363
R395 VSS.n49 VSS.n41 0.347226
R396 VSS.n67 VSS.n66 0.344944
R397 VSS.n71 VSS.n70 0.344944
R398 VSS.n43 VSS.n42 0.319807
R399 VSS.n46 VSS.n45 0.291342
R400 VSS.n49 VSS.n46 0.22669
R401 VSS.n77 VSS.n40 0.216409
R402 VSS.n130 VSS.n129 0.212
R403 VSS.n76 VSS.n54 0.210727
R404 VSS.n79 VSS.n78 0.158833
R405 VSS.n47 VSS.n46 0.158238
R406 VSS.n130 VSS 0.14
R407 VSS.n64 VSS.n59 0.135283
R408 VSS.n69 VSS.n57 0.135283
R409 VSS.n109 VSS.n108 0.120292
R410 VSS.n109 VSS.n104 0.120292
R411 VSS.n127 VSS.n105 0.120292
R412 VSS.n122 VSS.n105 0.120292
R413 VSS.n122 VSS.n121 0.120292
R414 VSS.n121 VSS.n116 0.120292
R415 VSS.n117 VSS.n116 0.120292
R416 VSS.n128 VSS.n104 0.112479
R417 VSS.n78 VSS.n77 0.09425
R418 VSS VSS.n132 0.0899516
R419 VSS.n45 VSS.n44 0.0714406
R420 VSS.n108 VSS 0.0603958
R421 VSS.n131 VSS.n0 0.0584812
R422 VSS VSS.n131 0.0520484
R423 VSS VSS.n1 0.0459545
R424 VSS.n102 VSS 0.0459545
R425 VSS.n68 VSS.n0 0.0455
R426 VSS.n33 VSS.n29 0.0429342
R427 VSS.n34 VSS.n33 0.0429342
R428 VSS.n35 VSS.n34 0.0429342
R429 VSS.n35 VSS.n28 0.0429342
R430 VSS.n31 VSS.n30 0.0389615
R431 VSS.n38 VSS.n28 0.0340526
R432 VSS.n1 VSS 0.0338333
R433 VSS.n102 VSS 0.0338333
R434 VSS.n46 VSS.n43 0.0289653
R435 VSS.n117 VSS 0.0226354
R436 VSS.n128 VSS.n127 0.0083125
R437 VSS.n31 VSS.n29 0.00773684
R438 VSS.n77 VSS.n76 0.00618182
R439 VSS.n131 VSS.n130 0.00544203
R440 VSS.n78 VSS.n0 0.00154167
R441 CTRL.n1 CTRL.t1 212.081
R442 CTRL.n25 CTRL.t3 212.081
R443 CTRL.n23 CTRL.t6 212.081
R444 CTRL.n2 CTRL.t12 212.081
R445 CTRL.n18 CTRL.t17 212.081
R446 CTRL.n3 CTRL.t0 212.081
R447 CTRL.n13 CTRL.t2 212.081
R448 CTRL.n11 CTRL.t4 212.081
R449 CTRL.n12 CTRL 163.264
R450 CTRL.n15 CTRL.n14 152
R451 CTRL.n17 CTRL.n16 152
R452 CTRL.n20 CTRL.n19 152
R453 CTRL.n22 CTRL.n21 152
R454 CTRL.n24 CTRL.n0 152
R455 CTRL CTRL.n26 152
R456 CTRL.n1 CTRL.t15 139.78
R457 CTRL.n25 CTRL.t11 139.78
R458 CTRL.n23 CTRL.t8 139.78
R459 CTRL.n2 CTRL.t10 139.78
R460 CTRL.n18 CTRL.t19 139.78
R461 CTRL.n3 CTRL.t5 139.78
R462 CTRL.n13 CTRL.t18 139.78
R463 CTRL.n11 CTRL.t13 139.78
R464 CTRL.n4 CTRL.t16 120.23
R465 CTRL.n4 CTRL.t9 120.228
R466 CTRL.n7 CTRL.t7 118.061
R467 CTRL.n7 CTRL.t14 118.058
R468 CTRL.n26 CTRL.n1 30.6732
R469 CTRL.n26 CTRL.n25 30.6732
R470 CTRL.n25 CTRL.n24 30.6732
R471 CTRL.n24 CTRL.n23 30.6732
R472 CTRL.n23 CTRL.n22 30.6732
R473 CTRL.n22 CTRL.n2 30.6732
R474 CTRL.n19 CTRL.n2 30.6732
R475 CTRL.n19 CTRL.n18 30.6732
R476 CTRL.n18 CTRL.n17 30.6732
R477 CTRL.n17 CTRL.n3 30.6732
R478 CTRL.n14 CTRL.n3 30.6732
R479 CTRL.n14 CTRL.n13 30.6732
R480 CTRL.n13 CTRL.n12 30.6732
R481 CTRL.n12 CTRL.n11 30.6732
R482 CTRL CTRL.n0 21.5045
R483 CTRL.n21 CTRL 19.4565
R484 CTRL CTRL.n20 17.4085
R485 CTRL CTRL.n15 13.3125
R486 CTRL.n16 CTRL.n10 13.0565
R487 CTRL.n15 CTRL 10.2405
R488 CTRL.n16 CTRL 8.1925
R489 CTRL.n20 CTRL 6.1445
R490 CTRL.n21 CTRL 4.0965
R491 CTRL.n10 CTRL.n9 3.2054
R492 CTRL.n10 CTRL 2.3045
R493 CTRL CTRL.n0 2.0485
R494 CTRL.n8 CTRL.n7 0.528909
R495 CTRL.n5 CTRL.n4 0.506182
R496 CTRL.n6 CTRL.n5 0.42675
R497 CTRL.n9 CTRL.n6 0.342556
R498 CTRL.n9 CTRL.n8 0.3415
R499 CTRL.n5 CTRL 0.170955
R500 CTRL.n8 CTRL 0.148227
R501 CTRL.n6 CTRL 0.01225
R502 OUT.n3 OUT.n1 199.941
R503 OUT.n10 OUT.n9 199.941
R504 OUT.n2 OUT.t7 83.7234
R505 OUT.n4 OUT.t6 83.7234
R506 OUT.n11 OUT.t0 83.7234
R507 OUT.n8 OUT.t1 83.7234
R508 OUT.n1 OUT.t2 28.5655
R509 OUT.n1 OUT.t3 28.5655
R510 OUT.n9 OUT.t5 28.5655
R511 OUT.n9 OUT.t4 28.5655
R512 OUT.n7 OUT.n6 1.15259
R513 OUT.n6 OUT.n5 0.938152
R514 OUT.n2 OUT.n0 0.5005
R515 OUT.n5 OUT.n4 0.5005
R516 OUT.n12 OUT.n11 0.5005
R517 OUT.n8 OUT.n7 0.5005
R518 OUT.n4 OUT.n3 0.478385
R519 OUT.n3 OUT.n2 0.478385
R520 OUT.n10 OUT.n8 0.478385
R521 OUT.n11 OUT.n10 0.478385
R522 OUT.n5 OUT.n0 0.364136
R523 OUT.n12 OUT.n7 0.364136
R524 OUT.n0 OUT 0.244818
R525 OUT OUT.n12 0.244818
R526 OUT.n6 OUT 0.0137188
C0 OUT myOpamp_0.INn 0.005273f
C1 a_1740_1605# tgate_1.IN 2.35765f
C2 IN a_1740_1605# 3.11184f
C3 sky130_fd_sc_hd__tap_2_0.VPB OUT 4.57e-19
C4 OUT VDD 2.99895f
C5 a_1998_1605# a_1740_1605# 1.57848f
C6 CTRL myOpamp_0.INn 0.25444f
C7 sky130_fd_sc_hd__tap_2_0.VPB CTRL 0.278876f
C8 a_944_1150# a_1740_1605# 0.27522f
C9 tgate_0.CTRL tgate_1.IN 1.18065f
C10 CTRL VDD 4.33897f
C11 IN tgate_0.CTRL 0.258603f
C12 myOpamp_0.INn a_1740_1605# 0.849481f
C13 a_1740_1605# VDD 4.48135f
C14 OUT CTRL 1.87653f
C15 myOpamp_0.INn tgate_0.CTRL 9.97e-19
C16 IN tgate_1.IN 0.820736f
C17 sky130_fd_sc_hd__tap_2_0.VPB tgate_0.CTRL 0.175567f
C18 a_1998_1605# tgate_1.IN 0.662032f
C19 tgate_0.CTRL VDD 4.18128f
C20 a_1998_1605# IN 0.763261f
C21 a_944_1150# tgate_1.IN 0.001336f
C22 a_944_1150# IN 0.197425f
C23 myOpamp_0.INn tgate_1.IN 1.8069f
C24 OUT tgate_0.CTRL 1.62697f
C25 IN myOpamp_0.INn 0.503808f
C26 a_944_1150# a_1998_1605# 1.5318f
C27 a_1998_1605# myOpamp_0.INn 1.23683f
C28 tgate_1.IN VDD 5.23603f
C29 IN VDD 6.85907f
C30 a_3626_n94# a_944_1150# 6.06e-20
C31 a_3626_n94# myOpamp_0.INn 0.007465f
C32 a_1998_1605# VDD 0.154599f
C33 CTRL tgate_0.CTRL 2.30483f
C34 a_944_1150# myOpamp_0.INn 1.1307f
C35 OUT tgate_1.IN 1.38344f
C36 OUT IN 1.3678f
C37 a_944_1150# VDD 0.125237f
C38 myOpamp_0.INn VDD 0.486138f
C39 sky130_fd_sc_hd__tap_2_0.VPB VDD 0.274328f
C40 CTRL tgate_1.IN 0.795971f
C41 CTRL IN 1.30918f
C42 OUT VSS 5.986641f
C43 IN VSS 11.177226f
C44 CTRL VSS 7.481905f
C45 VDD VSS 55.748493f
C46 tgate_0.CTRL VSS 4.58383f
C47 a_3626_n94# VSS 0.672562f
C48 a_944_1150# VSS 5.51409f
C49 a_1998_1605# VSS 1.65017f
C50 myOpamp_0.INn VSS 7.28783f
C51 tgate_1.IN VSS 2.60644f
C52 a_1740_1605# VSS 2.78479f
C53 sky130_fd_sc_hd__tap_2_0.VPB VSS 1.14309f
C54 OUT.n0 VSS 0.15064f
C55 OUT.t2 VSS 0.003712f
C56 OUT.t3 VSS 0.003712f
C57 OUT.n1 VSS 0.007689f
C58 OUT.t7 VSS 0.013418f
C59 OUT.n2 VSS 0.107926f
C60 OUT.n3 VSS 0.101076f
C61 OUT.t6 VSS 0.013275f
C62 OUT.n4 VSS 0.105508f
C63 OUT.n5 VSS 0.264386f
C64 OUT.n6 VSS 0.694965f
C65 OUT.n7 VSS 0.338431f
C66 OUT.t1 VSS 0.013275f
C67 OUT.n8 VSS 0.105508f
C68 OUT.t5 VSS 0.003712f
C69 OUT.t4 VSS 0.003712f
C70 OUT.n9 VSS 0.007689f
C71 OUT.n10 VSS 0.101076f
C72 OUT.t0 VSS 0.013418f
C73 OUT.n11 VSS 0.107926f
C74 OUT.n12 VSS 0.15064f
C75 CTRL.n0 VSS 0.005024f
C76 CTRL.t1 VSS 0.009174f
C77 CTRL.t15 VSS 0.005406f
C78 CTRL.n1 VSS 0.012365f
C79 CTRL.t3 VSS 0.009174f
C80 CTRL.t11 VSS 0.005406f
C81 CTRL.t6 VSS 0.009174f
C82 CTRL.t8 VSS 0.005406f
C83 CTRL.t12 VSS 0.009174f
C84 CTRL.t10 VSS 0.005406f
C85 CTRL.n2 VSS 0.01323f
C86 CTRL.t17 VSS 0.009174f
C87 CTRL.t19 VSS 0.005406f
C88 CTRL.t0 VSS 0.009174f
C89 CTRL.t5 VSS 0.005406f
C90 CTRL.n3 VSS 0.01323f
C91 CTRL.t16 VSS 0.102501f
C92 CTRL.t9 VSS 0.1025f
C93 CTRL.n4 VSS 0.565618f
C94 CTRL.n5 VSS 0.383326f
C95 CTRL.n6 VSS 1.06549f
C96 CTRL.t7 VSS 0.099823f
C97 CTRL.t14 VSS 0.099822f
C98 CTRL.n7 VSS 0.57775f
C99 CTRL.n8 VSS 0.379137f
C100 CTRL.n9 VSS 2.01491f
C101 CTRL.n10 VSS 0.308073f
C102 CTRL.t2 VSS 0.009174f
C103 CTRL.t18 VSS 0.005406f
C104 CTRL.t4 VSS 0.009174f
C105 CTRL.t13 VSS 0.005406f
C106 CTRL.n11 VSS 0.012365f
C107 CTRL.n12 VSS 0.006469f
C108 CTRL.n13 VSS 0.01323f
C109 CTRL.n14 VSS 0.006055f
C110 CTRL.n15 VSS 0.005024f
C111 CTRL.n16 VSS 0.004532f
C112 CTRL.n17 VSS 0.006055f
C113 CTRL.n18 VSS 0.01323f
C114 CTRL.n19 VSS 0.006055f
C115 CTRL.n20 VSS 0.005024f
C116 CTRL.n21 VSS 0.005024f
C117 CTRL.n22 VSS 0.006055f
C118 CTRL.n23 VSS 0.01323f
C119 CTRL.n24 VSS 0.006055f
C120 CTRL.n25 VSS 0.01323f
C121 CTRL.n26 VSS 0.006055f
C122 IN.t8 VSS 0.107729f
C123 IN.t6 VSS 0.107375f
C124 IN.n0 VSS 0.133f
C125 IN.t5 VSS 0.107375f
C126 IN.n1 VSS 0.078467f
C127 IN.t4 VSS 0.107375f
C128 IN.n2 VSS 0.068105f
C129 IN.t7 VSS 0.10765f
C130 IN.n3 VSS 0.18673f
C131 IN.t0 VSS 0.024658f
C132 IN.n4 VSS 0.095276f
C133 IN.t2 VSS 0.006818f
C134 IN.t1 VSS 0.006818f
C135 IN.n5 VSS 0.022125f
C136 IN.n6 VSS 0.134918f
C137 IN.t3 VSS 0.024658f
C138 IN.n7 VSS 0.071178f
C139 IN.n8 VSS 0.815587f
C140 IN.n9 VSS 3.13504f
C141 VDD.n0 VSS 0.684694f
C142 VDD.n1 VSS 0.741296f
C143 VDD.n2 VSS 0.121404f
C144 VDD.n3 VSS 0.121344f
C145 VDD.n4 VSS 0.242837f
C146 VDD.n5 VSS 0.243017f
C147 VDD.n6 VSS 0.738083f
C148 VDD.n7 VSS 0.121284f
C149 VDD.n8 VSS 0.121674f
C150 VDD.n9 VSS 0.725268f
C151 VDD.n10 VSS 0.120961f
C152 VDD.n11 VSS 0.120575f
C153 VDD.n12 VSS 0.241386f
C154 VDD.n13 VSS 0.724332f
C155 VDD.n14 VSS 0.740837f
C156 VDD.n15 VSS 0.726204f
C157 VDD.n16 VSS 0.241628f
C158 VDD.n17 VSS 0.120783f
C159 VDD.n18 VSS 0.120843f
C160 VDD.n19 VSS 0.415513f
C161 VDD.n20 VSS 0.775247f
C162 VDD.t10 VSS 0.04254f
C163 VDD.t12 VSS 0.009634f
C164 VDD.n21 VSS 0.055744f
C165 VDD.t21 VSS 0.002622f
C166 VDD.t27 VSS 0.002622f
C167 VDD.n22 VSS 0.005422f
C168 VDD.n23 VSS 0.107667f
C169 VDD.t35 VSS 0.002622f
C170 VDD.t33 VSS 0.002622f
C171 VDD.n24 VSS 0.005422f
C172 VDD.n25 VSS 0.090512f
C173 VDD.t13 VSS 0.042512f
C174 VDD.t15 VSS 0.009634f
C175 VDD.n26 VSS 0.096515f
C176 VDD.t23 VSS 0.002622f
C177 VDD.t29 VSS 0.002622f
C178 VDD.n27 VSS 0.005422f
C179 VDD.n28 VSS 0.12928f
C180 VDD.t19 VSS 0.002622f
C181 VDD.t25 VSS 0.002622f
C182 VDD.n29 VSS 0.005422f
C183 VDD.n30 VSS 0.07912f
C184 VDD.t11 VSS 0.149525f
C185 VDD.t20 VSS 0.119435f
C186 VDD.t26 VSS 0.119435f
C187 VDD.t34 VSS 0.119435f
C188 VDD.t32 VSS 0.119435f
C189 VDD.t30 VSS 0.085873f
C190 VDD.t14 VSS 0.149525f
C191 VDD.t28 VSS 0.119435f
C192 VDD.t22 VSS 0.119435f
C193 VDD.t24 VSS 0.119435f
C194 VDD.t18 VSS 0.119435f
C195 VDD.t16 VSS 0.09328f
C196 VDD.n31 VSS -0.07004f
C197 VDD.t8 VSS 0.098222f
C198 VDD.n32 VSS 0.151915f
C199 VDD.n33 VSS 0.020615f
C200 VDD.t31 VSS 0.002622f
C201 VDD.t17 VSS 0.002622f
C202 VDD.n34 VSS 0.005422f
C203 VDD.n35 VSS 0.088966f
C204 VDD.n36 VSS 3.16909f
C205 VDD.n37 VSS 0.031918f
C206 VDD.n38 VSS 0.018396f
C207 VDD.n39 VSS 0.131297f
C208 VDD.t7 VSS 0.104678f
C209 VDD.n40 VSS 0.066249f
C210 VDD.t0 VSS 0.104678f
C211 VDD.n41 VSS 0.108462f
C212 VDD.n42 VSS 0.056763f
C213 VDD.n43 VSS 0.250093f
C214 VDD.n44 VSS 0.031918f
C215 VDD.n45 VSS 0.018396f
C216 VDD.n46 VSS 0.131297f
C217 VDD.t5 VSS 0.104678f
C218 VDD.n47 VSS 0.066249f
C219 VDD.t6 VSS 0.104678f
C220 VDD.n48 VSS 0.108462f
C221 VDD.n49 VSS 0.056763f
C222 VDD.n50 VSS 0.253193f
C223 VDD.n51 VSS 0.423703f
C224 VDD.n52 VSS 0.004166f
C225 VDD.n53 VSS 0.007985f
C226 VDD.t3 VSS 0.002441f
C227 VDD.t4 VSS 0.002441f
C228 VDD.n54 VSS 0.00524f
C229 VDD.t2 VSS 0.002441f
C230 VDD.t37 VSS 0.002441f
C231 VDD.n55 VSS 0.00524f
C232 VDD.n56 VSS 0.002183f
C233 VDD.t9 VSS 0.009294f
C234 VDD.n57 VSS 0.013242f
C235 VDD.n58 VSS 0.005989f
C236 VDD.n59 VSS 0.007985f
C237 VDD.n60 VSS 0.007985f
C238 VDD.n61 VSS 0.001552f
C239 VDD.n62 VSS 0.005975f
C240 VDD.n63 VSS 0.002582f
C241 VDD.n64 VSS 0.005975f
C242 VDD.t38 VSS 0.002441f
C243 VDD.t36 VSS 0.002441f
C244 VDD.n65 VSS 0.00524f
C245 VDD.n66 VSS 0.001967f
C246 VDD.t1 VSS 0.009295f
C247 VDD.n67 VSS 0.010924f
C248 VDD.n68 VSS 0.004982f
C249 VDD.n69 VSS 0.007985f
C250 VDD.n70 VSS 0.007985f
C251 VDD.n71 VSS 0.001768f
C252 VDD.n72 VSS 0.005975f
C253 VDD.n73 VSS 0.002475f
C254 VDD.n74 VSS 0.001522f
C255 VDD.n75 VSS 0.007812f
C256 VDD.n76 VSS 0.320945f
C257 VDD.n77 VSS 4.09192f
C258 VDD.n78 VSS 2.91201f
C259 VDD.n79 VSS 1.55711f
C260 VDD.n80 VSS 0.730917f
.ends

