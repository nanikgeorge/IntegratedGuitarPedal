magic
tech sky130A
magscale 1 2
timestamp 1713312949
<< nmos >>
rect -100 -469 100 531
<< ndiff >>
rect -158 519 -100 531
rect -158 -457 -146 519
rect -112 -457 -100 519
rect -158 -469 -100 -457
rect 100 519 158 531
rect 100 -457 112 519
rect 146 -457 158 519
rect 100 -469 158 -457
<< ndiffc >>
rect -146 -457 -112 519
rect 112 -457 146 519
<< poly >>
rect -100 531 100 557
rect -100 -507 100 -469
rect -100 -541 -84 -507
rect 84 -541 100 -507
rect -100 -557 100 -541
<< polycont >>
rect -84 -541 84 -507
<< locali >>
rect -146 519 -112 535
rect -146 -473 -112 -457
rect 112 519 146 535
rect 112 -473 146 -457
rect -100 -541 -84 -507
rect 84 -541 100 -507
<< viali >>
rect -146 -457 -112 519
rect 112 -457 146 519
rect -84 -541 84 -507
<< metal1 >>
rect -152 519 -106 531
rect -152 -457 -146 519
rect -112 -457 -106 519
rect -152 -469 -106 -457
rect 106 519 152 531
rect 106 -457 112 519
rect 146 -457 152 519
rect 106 -469 152 -457
rect -96 -507 96 -501
rect -96 -541 -84 -507
rect 84 -541 96 -507
rect -96 -547 96 -541
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5 l 1 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
