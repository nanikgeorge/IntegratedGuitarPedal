magic
tech sky130A
magscale 1 2
timestamp 1713533072
<< nwell >>
rect 5616 37798 11316 37998
rect 5616 35398 5816 37798
rect 7442 36810 10668 37322
rect 11116 35398 11316 37798
rect 12723 37963 13573 38531
rect 18404 37916 24104 38116
rect 12723 36503 13573 37071
rect 18404 35516 18604 37916
rect 20230 36928 23456 37440
rect 23904 35516 24104 37916
rect 25511 38081 26361 38649
rect 5616 35198 11316 35398
rect 12516 35167 13604 35488
rect 18404 35316 24104 35516
rect 25511 36621 26361 37189
rect 25304 35285 26392 35606
rect 5636 31872 11336 32072
rect 5636 29472 5836 31872
rect 7462 30884 10688 31396
rect 11136 29472 11336 31872
rect 12743 32037 13593 32605
rect 5636 29272 11336 29472
rect 18368 31796 24068 31996
rect 12743 30577 13593 31145
rect 12536 29241 13624 29562
rect 18368 29396 18568 31796
rect 20194 30808 23420 31320
rect 23868 29396 24068 31796
rect 25475 31961 26325 32529
rect 18368 29196 24068 29396
rect 25475 30501 26325 31069
rect 25268 29165 26356 29486
rect 5756 25168 11456 25368
rect 5756 22768 5956 25168
rect 7582 24180 10808 24692
rect 11256 22768 11456 25168
rect 12863 25333 13713 25901
rect 5756 22568 11456 22768
rect 18464 25038 24164 25238
rect 12863 23873 13713 24441
rect 12656 22537 13744 22858
rect 18464 22638 18664 25038
rect 20290 24050 23516 24562
rect 23964 22638 24164 25038
rect 25571 25203 26421 25771
rect 18464 22438 24164 22638
rect 25571 23743 26421 24311
rect 25364 22407 26452 22728
rect 5632 18122 11332 18322
rect 5632 15722 5832 18122
rect 7458 17134 10684 17646
rect 11132 15722 11332 18122
rect 12739 18287 13589 18855
rect 5632 15522 11332 15722
rect 18814 17992 24514 18192
rect 12739 16827 13589 17395
rect 12532 15491 13620 15812
rect 18814 15592 19014 17992
rect 20640 17004 23866 17516
rect 24314 15592 24514 17992
rect 25921 18157 26771 18725
rect 18814 15392 24514 15592
rect 25921 16697 26771 17265
rect 25714 15361 26802 15682
<< pwell >>
rect 5916 37498 11016 37698
rect 5916 35698 7406 37498
rect 7436 35928 10666 36098
rect 10816 35698 11016 37498
rect 5916 35498 11016 35698
rect 12723 37405 13573 37963
rect 12723 35945 13573 36503
rect 18704 37616 23804 37816
rect 18704 35816 20194 37616
rect 20224 36046 23454 36216
rect 23604 35816 23804 37616
rect 18704 35616 23804 35816
rect 12588 34927 13362 35109
rect 13385 34944 13563 35101
rect 12588 34923 12617 34927
rect 12583 34889 12617 34923
rect 22244 34736 24208 35206
rect 24244 34736 24714 37900
rect 25511 37523 26361 38081
rect 25511 36063 26361 36621
rect 25376 35045 26150 35227
rect 26173 35062 26351 35219
rect 25376 35041 25405 35045
rect 25371 35007 25405 35041
rect 5936 31572 11036 31772
rect 5936 29772 7426 31572
rect 7456 30002 10686 30172
rect 10836 29772 11036 31572
rect 5936 29572 11036 29772
rect 9476 28692 11440 29162
rect 11476 28692 11946 31856
rect 12743 31479 13593 32037
rect 12743 30019 13593 30577
rect 18668 31496 23768 31696
rect 18668 29696 20158 31496
rect 20188 29926 23418 30096
rect 23568 29696 23768 31496
rect 18668 29496 23768 29696
rect 12608 29001 13382 29183
rect 13405 29018 13583 29175
rect 12608 28997 12637 29001
rect 12603 28963 12637 28997
rect 22208 28616 24172 29086
rect 24208 28616 24678 31780
rect 25475 31403 26325 31961
rect 25475 29943 26325 30501
rect 25340 28925 26114 29107
rect 26137 28942 26315 29099
rect 25340 28921 25369 28925
rect 25335 28887 25369 28921
rect 6056 24868 11156 25068
rect 6056 23068 7546 24868
rect 7576 23298 10806 23468
rect 10956 23068 11156 24868
rect 6056 22868 11156 23068
rect 9596 21988 11560 22458
rect 11596 21988 12066 25152
rect 12863 24775 13713 25333
rect 12863 23315 13713 23873
rect 18764 24738 23864 24938
rect 18764 22938 20254 24738
rect 20284 23168 23514 23338
rect 23664 22938 23864 24738
rect 18764 22738 23864 22938
rect 12728 22297 13502 22479
rect 13525 22314 13703 22471
rect 12728 22293 12757 22297
rect 12723 22259 12757 22293
rect 22304 21858 24268 22328
rect 24304 21858 24774 25022
rect 25571 24645 26421 25203
rect 25571 23185 26421 23743
rect 25436 22167 26210 22349
rect 26233 22184 26411 22341
rect 25436 22163 25465 22167
rect 25431 22129 25465 22163
rect 5932 17822 11032 18022
rect 5932 16022 7422 17822
rect 7452 16252 10682 16422
rect 10832 16022 11032 17822
rect 5932 15822 11032 16022
rect 9472 14942 11436 15412
rect 11472 14942 11942 18106
rect 12739 17729 13589 18287
rect 12739 16269 13589 16827
rect 19114 17692 24214 17892
rect 19114 15892 20604 17692
rect 20634 16122 23864 16292
rect 24014 15892 24214 17692
rect 19114 15692 24214 15892
rect 12604 15251 13378 15433
rect 13401 15268 13579 15425
rect 12604 15247 12633 15251
rect 12599 15213 12633 15247
rect 22654 14812 24618 15282
rect 24654 14812 25124 17976
rect 25921 17599 26771 18157
rect 25921 16139 26771 16697
rect 25786 15121 26560 15303
rect 26583 15138 26761 15295
rect 25786 15117 25815 15121
rect 25781 15083 25815 15117
<< nmos >>
rect 7536 36483 7736 36683
rect 7794 36483 7994 36683
rect 8052 36483 8252 36683
rect 8310 36483 8510 36683
rect 8568 36483 8768 36683
rect 8826 36483 9026 36683
rect 9084 36483 9284 36683
rect 9342 36483 9542 36683
rect 9600 36483 9800 36683
rect 9858 36483 10058 36683
rect 10116 36483 10316 36683
rect 10374 36483 10574 36683
rect 7536 36163 7736 36247
rect 7794 36163 7994 36247
rect 8052 36163 8252 36247
rect 8310 36163 8510 36247
rect 8568 36163 8768 36247
rect 8826 36163 9026 36247
rect 9084 36163 9284 36247
rect 9342 36163 9542 36247
rect 9600 36163 9800 36247
rect 9858 36163 10058 36247
rect 10116 36163 10316 36247
rect 10374 36163 10574 36247
rect 12919 37615 13119 37815
rect 13177 37615 13377 37815
rect 12919 36155 13119 36355
rect 13177 36155 13377 36355
rect 20324 36601 20524 36801
rect 20582 36601 20782 36801
rect 20840 36601 21040 36801
rect 21098 36601 21298 36801
rect 21356 36601 21556 36801
rect 21614 36601 21814 36801
rect 21872 36601 22072 36801
rect 22130 36601 22330 36801
rect 22388 36601 22588 36801
rect 22646 36601 22846 36801
rect 22904 36601 23104 36801
rect 23162 36601 23362 36801
rect 20324 36281 20524 36365
rect 20582 36281 20782 36365
rect 20840 36281 21040 36365
rect 21098 36281 21298 36365
rect 21356 36281 21556 36365
rect 21614 36281 21814 36365
rect 21872 36281 22072 36365
rect 22130 36281 22330 36365
rect 22388 36281 22588 36365
rect 22646 36281 22846 36365
rect 22904 36281 23104 36365
rect 23162 36281 23362 36365
rect 25707 37733 25907 37933
rect 25965 37733 26165 37933
rect 25707 36273 25907 36473
rect 25965 36273 26165 36473
rect 7556 30557 7756 30757
rect 7814 30557 8014 30757
rect 8072 30557 8272 30757
rect 8330 30557 8530 30757
rect 8588 30557 8788 30757
rect 8846 30557 9046 30757
rect 9104 30557 9304 30757
rect 9362 30557 9562 30757
rect 9620 30557 9820 30757
rect 9878 30557 10078 30757
rect 10136 30557 10336 30757
rect 10394 30557 10594 30757
rect 7556 30237 7756 30321
rect 7814 30237 8014 30321
rect 8072 30237 8272 30321
rect 8330 30237 8530 30321
rect 8588 30237 8788 30321
rect 8846 30237 9046 30321
rect 9104 30237 9304 30321
rect 9362 30237 9562 30321
rect 9620 30237 9820 30321
rect 9878 30237 10078 30321
rect 10136 30237 10336 30321
rect 10394 30237 10594 30321
rect 12939 31689 13139 31889
rect 13197 31689 13397 31889
rect 12939 30229 13139 30429
rect 13197 30229 13397 30429
rect 20288 30481 20488 30681
rect 20546 30481 20746 30681
rect 20804 30481 21004 30681
rect 21062 30481 21262 30681
rect 21320 30481 21520 30681
rect 21578 30481 21778 30681
rect 21836 30481 22036 30681
rect 22094 30481 22294 30681
rect 22352 30481 22552 30681
rect 22610 30481 22810 30681
rect 22868 30481 23068 30681
rect 23126 30481 23326 30681
rect 20288 30161 20488 30245
rect 20546 30161 20746 30245
rect 20804 30161 21004 30245
rect 21062 30161 21262 30245
rect 21320 30161 21520 30245
rect 21578 30161 21778 30245
rect 21836 30161 22036 30245
rect 22094 30161 22294 30245
rect 22352 30161 22552 30245
rect 22610 30161 22810 30245
rect 22868 30161 23068 30245
rect 23126 30161 23326 30245
rect 25671 31613 25871 31813
rect 25929 31613 26129 31813
rect 25671 30153 25871 30353
rect 25929 30153 26129 30353
rect 7676 23853 7876 24053
rect 7934 23853 8134 24053
rect 8192 23853 8392 24053
rect 8450 23853 8650 24053
rect 8708 23853 8908 24053
rect 8966 23853 9166 24053
rect 9224 23853 9424 24053
rect 9482 23853 9682 24053
rect 9740 23853 9940 24053
rect 9998 23853 10198 24053
rect 10256 23853 10456 24053
rect 10514 23853 10714 24053
rect 7676 23533 7876 23617
rect 7934 23533 8134 23617
rect 8192 23533 8392 23617
rect 8450 23533 8650 23617
rect 8708 23533 8908 23617
rect 8966 23533 9166 23617
rect 9224 23533 9424 23617
rect 9482 23533 9682 23617
rect 9740 23533 9940 23617
rect 9998 23533 10198 23617
rect 10256 23533 10456 23617
rect 10514 23533 10714 23617
rect 13059 24985 13259 25185
rect 13317 24985 13517 25185
rect 13059 23525 13259 23725
rect 13317 23525 13517 23725
rect 20384 23723 20584 23923
rect 20642 23723 20842 23923
rect 20900 23723 21100 23923
rect 21158 23723 21358 23923
rect 21416 23723 21616 23923
rect 21674 23723 21874 23923
rect 21932 23723 22132 23923
rect 22190 23723 22390 23923
rect 22448 23723 22648 23923
rect 22706 23723 22906 23923
rect 22964 23723 23164 23923
rect 23222 23723 23422 23923
rect 20384 23403 20584 23487
rect 20642 23403 20842 23487
rect 20900 23403 21100 23487
rect 21158 23403 21358 23487
rect 21416 23403 21616 23487
rect 21674 23403 21874 23487
rect 21932 23403 22132 23487
rect 22190 23403 22390 23487
rect 22448 23403 22648 23487
rect 22706 23403 22906 23487
rect 22964 23403 23164 23487
rect 23222 23403 23422 23487
rect 25767 24855 25967 25055
rect 26025 24855 26225 25055
rect 25767 23395 25967 23595
rect 26025 23395 26225 23595
rect 7552 16807 7752 17007
rect 7810 16807 8010 17007
rect 8068 16807 8268 17007
rect 8326 16807 8526 17007
rect 8584 16807 8784 17007
rect 8842 16807 9042 17007
rect 9100 16807 9300 17007
rect 9358 16807 9558 17007
rect 9616 16807 9816 17007
rect 9874 16807 10074 17007
rect 10132 16807 10332 17007
rect 10390 16807 10590 17007
rect 7552 16487 7752 16571
rect 7810 16487 8010 16571
rect 8068 16487 8268 16571
rect 8326 16487 8526 16571
rect 8584 16487 8784 16571
rect 8842 16487 9042 16571
rect 9100 16487 9300 16571
rect 9358 16487 9558 16571
rect 9616 16487 9816 16571
rect 9874 16487 10074 16571
rect 10132 16487 10332 16571
rect 10390 16487 10590 16571
rect 12935 17939 13135 18139
rect 13193 17939 13393 18139
rect 12935 16479 13135 16679
rect 13193 16479 13393 16679
rect 20734 16677 20934 16877
rect 20992 16677 21192 16877
rect 21250 16677 21450 16877
rect 21508 16677 21708 16877
rect 21766 16677 21966 16877
rect 22024 16677 22224 16877
rect 22282 16677 22482 16877
rect 22540 16677 22740 16877
rect 22798 16677 22998 16877
rect 23056 16677 23256 16877
rect 23314 16677 23514 16877
rect 23572 16677 23772 16877
rect 20734 16357 20934 16441
rect 20992 16357 21192 16441
rect 21250 16357 21450 16441
rect 21508 16357 21708 16441
rect 21766 16357 21966 16441
rect 22024 16357 22224 16441
rect 22282 16357 22482 16441
rect 22540 16357 22740 16441
rect 22798 16357 22998 16441
rect 23056 16357 23256 16441
rect 23314 16357 23514 16441
rect 23572 16357 23772 16441
rect 26117 17809 26317 18009
rect 26375 17809 26575 18009
rect 26117 16349 26317 16549
rect 26375 16349 26575 16549
<< scnmos >>
rect 12666 34953 12696 35083
rect 12750 34953 12780 35083
rect 12834 34953 12864 35083
rect 12918 34953 12948 35083
rect 13002 34953 13032 35083
rect 13086 34953 13116 35083
rect 13170 34953 13200 35083
rect 13254 34953 13284 35083
rect 25454 35071 25484 35201
rect 25538 35071 25568 35201
rect 25622 35071 25652 35201
rect 25706 35071 25736 35201
rect 25790 35071 25820 35201
rect 25874 35071 25904 35201
rect 25958 35071 25988 35201
rect 26042 35071 26072 35201
rect 12686 29027 12716 29157
rect 12770 29027 12800 29157
rect 12854 29027 12884 29157
rect 12938 29027 12968 29157
rect 13022 29027 13052 29157
rect 13106 29027 13136 29157
rect 13190 29027 13220 29157
rect 13274 29027 13304 29157
rect 25418 28951 25448 29081
rect 25502 28951 25532 29081
rect 25586 28951 25616 29081
rect 25670 28951 25700 29081
rect 25754 28951 25784 29081
rect 25838 28951 25868 29081
rect 25922 28951 25952 29081
rect 26006 28951 26036 29081
rect 12806 22323 12836 22453
rect 12890 22323 12920 22453
rect 12974 22323 13004 22453
rect 13058 22323 13088 22453
rect 13142 22323 13172 22453
rect 13226 22323 13256 22453
rect 13310 22323 13340 22453
rect 13394 22323 13424 22453
rect 25514 22193 25544 22323
rect 25598 22193 25628 22323
rect 25682 22193 25712 22323
rect 25766 22193 25796 22323
rect 25850 22193 25880 22323
rect 25934 22193 25964 22323
rect 26018 22193 26048 22323
rect 26102 22193 26132 22323
rect 12682 15277 12712 15407
rect 12766 15277 12796 15407
rect 12850 15277 12880 15407
rect 12934 15277 12964 15407
rect 13018 15277 13048 15407
rect 13102 15277 13132 15407
rect 13186 15277 13216 15407
rect 13270 15277 13300 15407
rect 25864 15147 25894 15277
rect 25948 15147 25978 15277
rect 26032 15147 26062 15277
rect 26116 15147 26146 15277
rect 26200 15147 26230 15277
rect 26284 15147 26314 15277
rect 26368 15147 26398 15277
rect 26452 15147 26482 15277
<< pmos >>
rect 12919 38111 13119 38311
rect 13177 38111 13377 38311
rect 25707 38229 25907 38429
rect 25965 38229 26165 38429
rect 7536 36910 7736 37110
rect 7794 36910 7994 37110
rect 8052 36910 8252 37110
rect 8310 36910 8510 37110
rect 8568 36910 8768 37110
rect 8826 36910 9026 37110
rect 9084 36910 9284 37110
rect 9342 36910 9542 37110
rect 9600 36910 9800 37110
rect 9858 36910 10058 37110
rect 10116 36910 10316 37110
rect 10374 36910 10574 37110
rect 12919 36651 13119 36851
rect 13177 36651 13377 36851
rect 20324 37028 20524 37228
rect 20582 37028 20782 37228
rect 20840 37028 21040 37228
rect 21098 37028 21298 37228
rect 21356 37028 21556 37228
rect 21614 37028 21814 37228
rect 21872 37028 22072 37228
rect 22130 37028 22330 37228
rect 22388 37028 22588 37228
rect 22646 37028 22846 37228
rect 22904 37028 23104 37228
rect 23162 37028 23362 37228
rect 25707 36769 25907 36969
rect 25965 36769 26165 36969
rect 12939 32185 13139 32385
rect 13197 32185 13397 32385
rect 25671 32109 25871 32309
rect 25929 32109 26129 32309
rect 7556 30984 7756 31184
rect 7814 30984 8014 31184
rect 8072 30984 8272 31184
rect 8330 30984 8530 31184
rect 8588 30984 8788 31184
rect 8846 30984 9046 31184
rect 9104 30984 9304 31184
rect 9362 30984 9562 31184
rect 9620 30984 9820 31184
rect 9878 30984 10078 31184
rect 10136 30984 10336 31184
rect 10394 30984 10594 31184
rect 12939 30725 13139 30925
rect 13197 30725 13397 30925
rect 20288 30908 20488 31108
rect 20546 30908 20746 31108
rect 20804 30908 21004 31108
rect 21062 30908 21262 31108
rect 21320 30908 21520 31108
rect 21578 30908 21778 31108
rect 21836 30908 22036 31108
rect 22094 30908 22294 31108
rect 22352 30908 22552 31108
rect 22610 30908 22810 31108
rect 22868 30908 23068 31108
rect 23126 30908 23326 31108
rect 25671 30649 25871 30849
rect 25929 30649 26129 30849
rect 13059 25481 13259 25681
rect 13317 25481 13517 25681
rect 25767 25351 25967 25551
rect 26025 25351 26225 25551
rect 7676 24280 7876 24480
rect 7934 24280 8134 24480
rect 8192 24280 8392 24480
rect 8450 24280 8650 24480
rect 8708 24280 8908 24480
rect 8966 24280 9166 24480
rect 9224 24280 9424 24480
rect 9482 24280 9682 24480
rect 9740 24280 9940 24480
rect 9998 24280 10198 24480
rect 10256 24280 10456 24480
rect 10514 24280 10714 24480
rect 13059 24021 13259 24221
rect 13317 24021 13517 24221
rect 20384 24150 20584 24350
rect 20642 24150 20842 24350
rect 20900 24150 21100 24350
rect 21158 24150 21358 24350
rect 21416 24150 21616 24350
rect 21674 24150 21874 24350
rect 21932 24150 22132 24350
rect 22190 24150 22390 24350
rect 22448 24150 22648 24350
rect 22706 24150 22906 24350
rect 22964 24150 23164 24350
rect 23222 24150 23422 24350
rect 25767 23891 25967 24091
rect 26025 23891 26225 24091
rect 12935 18435 13135 18635
rect 13193 18435 13393 18635
rect 26117 18305 26317 18505
rect 26375 18305 26575 18505
rect 7552 17234 7752 17434
rect 7810 17234 8010 17434
rect 8068 17234 8268 17434
rect 8326 17234 8526 17434
rect 8584 17234 8784 17434
rect 8842 17234 9042 17434
rect 9100 17234 9300 17434
rect 9358 17234 9558 17434
rect 9616 17234 9816 17434
rect 9874 17234 10074 17434
rect 10132 17234 10332 17434
rect 10390 17234 10590 17434
rect 12935 16975 13135 17175
rect 13193 16975 13393 17175
rect 20734 17104 20934 17304
rect 20992 17104 21192 17304
rect 21250 17104 21450 17304
rect 21508 17104 21708 17304
rect 21766 17104 21966 17304
rect 22024 17104 22224 17304
rect 22282 17104 22482 17304
rect 22540 17104 22740 17304
rect 22798 17104 22998 17304
rect 23056 17104 23256 17304
rect 23314 17104 23514 17304
rect 23572 17104 23772 17304
rect 26117 16845 26317 17045
rect 26375 16845 26575 17045
<< scpmoshvt >>
rect 12666 35203 12696 35403
rect 12750 35203 12780 35403
rect 12834 35203 12864 35403
rect 12918 35203 12948 35403
rect 13002 35203 13032 35403
rect 13086 35203 13116 35403
rect 13170 35203 13200 35403
rect 13254 35203 13284 35403
rect 25454 35321 25484 35521
rect 25538 35321 25568 35521
rect 25622 35321 25652 35521
rect 25706 35321 25736 35521
rect 25790 35321 25820 35521
rect 25874 35321 25904 35521
rect 25958 35321 25988 35521
rect 26042 35321 26072 35521
rect 12686 29277 12716 29477
rect 12770 29277 12800 29477
rect 12854 29277 12884 29477
rect 12938 29277 12968 29477
rect 13022 29277 13052 29477
rect 13106 29277 13136 29477
rect 13190 29277 13220 29477
rect 13274 29277 13304 29477
rect 25418 29201 25448 29401
rect 25502 29201 25532 29401
rect 25586 29201 25616 29401
rect 25670 29201 25700 29401
rect 25754 29201 25784 29401
rect 25838 29201 25868 29401
rect 25922 29201 25952 29401
rect 26006 29201 26036 29401
rect 12806 22573 12836 22773
rect 12890 22573 12920 22773
rect 12974 22573 13004 22773
rect 13058 22573 13088 22773
rect 13142 22573 13172 22773
rect 13226 22573 13256 22773
rect 13310 22573 13340 22773
rect 13394 22573 13424 22773
rect 25514 22443 25544 22643
rect 25598 22443 25628 22643
rect 25682 22443 25712 22643
rect 25766 22443 25796 22643
rect 25850 22443 25880 22643
rect 25934 22443 25964 22643
rect 26018 22443 26048 22643
rect 26102 22443 26132 22643
rect 12682 15527 12712 15727
rect 12766 15527 12796 15727
rect 12850 15527 12880 15727
rect 12934 15527 12964 15727
rect 13018 15527 13048 15727
rect 13102 15527 13132 15727
rect 13186 15527 13216 15727
rect 13270 15527 13300 15727
rect 25864 15397 25894 15597
rect 25948 15397 25978 15597
rect 26032 15397 26062 15597
rect 26116 15397 26146 15597
rect 26200 15397 26230 15597
rect 26284 15397 26314 15597
rect 26368 15397 26398 15597
rect 26452 15397 26482 15597
<< ndiff >>
rect 7478 36671 7536 36683
rect 7478 36495 7490 36671
rect 7524 36495 7536 36671
rect 7478 36483 7536 36495
rect 7736 36671 7794 36683
rect 7736 36495 7748 36671
rect 7782 36495 7794 36671
rect 7736 36483 7794 36495
rect 7994 36671 8052 36683
rect 7994 36495 8006 36671
rect 8040 36495 8052 36671
rect 7994 36483 8052 36495
rect 8252 36671 8310 36683
rect 8252 36495 8264 36671
rect 8298 36495 8310 36671
rect 8252 36483 8310 36495
rect 8510 36671 8568 36683
rect 8510 36495 8522 36671
rect 8556 36495 8568 36671
rect 8510 36483 8568 36495
rect 8768 36671 8826 36683
rect 8768 36495 8780 36671
rect 8814 36495 8826 36671
rect 8768 36483 8826 36495
rect 9026 36671 9084 36683
rect 9026 36495 9038 36671
rect 9072 36495 9084 36671
rect 9026 36483 9084 36495
rect 9284 36671 9342 36683
rect 9284 36495 9296 36671
rect 9330 36495 9342 36671
rect 9284 36483 9342 36495
rect 9542 36671 9600 36683
rect 9542 36495 9554 36671
rect 9588 36495 9600 36671
rect 9542 36483 9600 36495
rect 9800 36671 9858 36683
rect 9800 36495 9812 36671
rect 9846 36495 9858 36671
rect 9800 36483 9858 36495
rect 10058 36671 10116 36683
rect 10058 36495 10070 36671
rect 10104 36495 10116 36671
rect 10058 36483 10116 36495
rect 10316 36671 10374 36683
rect 10316 36495 10328 36671
rect 10362 36495 10374 36671
rect 10316 36483 10374 36495
rect 10574 36671 10632 36683
rect 10574 36495 10586 36671
rect 10620 36495 10632 36671
rect 10574 36483 10632 36495
rect 7478 36235 7536 36247
rect 7478 36175 7490 36235
rect 7524 36175 7536 36235
rect 7478 36163 7536 36175
rect 7736 36235 7794 36247
rect 7736 36175 7748 36235
rect 7782 36175 7794 36235
rect 7736 36163 7794 36175
rect 7994 36235 8052 36247
rect 7994 36175 8006 36235
rect 8040 36175 8052 36235
rect 7994 36163 8052 36175
rect 8252 36235 8310 36247
rect 8252 36175 8264 36235
rect 8298 36175 8310 36235
rect 8252 36163 8310 36175
rect 8510 36235 8568 36247
rect 8510 36175 8522 36235
rect 8556 36175 8568 36235
rect 8510 36163 8568 36175
rect 8768 36235 8826 36247
rect 8768 36175 8780 36235
rect 8814 36175 8826 36235
rect 8768 36163 8826 36175
rect 9026 36235 9084 36247
rect 9026 36175 9038 36235
rect 9072 36175 9084 36235
rect 9026 36163 9084 36175
rect 9284 36235 9342 36247
rect 9284 36175 9296 36235
rect 9330 36175 9342 36235
rect 9284 36163 9342 36175
rect 9542 36235 9600 36247
rect 9542 36175 9554 36235
rect 9588 36175 9600 36235
rect 9542 36163 9600 36175
rect 9800 36235 9858 36247
rect 9800 36175 9812 36235
rect 9846 36175 9858 36235
rect 9800 36163 9858 36175
rect 10058 36235 10116 36247
rect 10058 36175 10070 36235
rect 10104 36175 10116 36235
rect 10058 36163 10116 36175
rect 10316 36235 10374 36247
rect 10316 36175 10328 36235
rect 10362 36175 10374 36235
rect 10316 36163 10374 36175
rect 10574 36235 10632 36247
rect 10574 36175 10586 36235
rect 10620 36175 10632 36235
rect 10574 36163 10632 36175
rect 12861 37803 12919 37815
rect 12861 37627 12873 37803
rect 12907 37627 12919 37803
rect 12861 37615 12919 37627
rect 13119 37803 13177 37815
rect 13119 37627 13131 37803
rect 13165 37627 13177 37803
rect 13119 37615 13177 37627
rect 13377 37803 13435 37815
rect 13377 37627 13389 37803
rect 13423 37627 13435 37803
rect 13377 37615 13435 37627
rect 12861 36343 12919 36355
rect 12861 36167 12873 36343
rect 12907 36167 12919 36343
rect 12861 36155 12919 36167
rect 13119 36343 13177 36355
rect 13119 36167 13131 36343
rect 13165 36167 13177 36343
rect 13119 36155 13177 36167
rect 13377 36343 13435 36355
rect 13377 36167 13389 36343
rect 13423 36167 13435 36343
rect 13377 36155 13435 36167
rect 20266 36789 20324 36801
rect 20266 36613 20278 36789
rect 20312 36613 20324 36789
rect 20266 36601 20324 36613
rect 20524 36789 20582 36801
rect 20524 36613 20536 36789
rect 20570 36613 20582 36789
rect 20524 36601 20582 36613
rect 20782 36789 20840 36801
rect 20782 36613 20794 36789
rect 20828 36613 20840 36789
rect 20782 36601 20840 36613
rect 21040 36789 21098 36801
rect 21040 36613 21052 36789
rect 21086 36613 21098 36789
rect 21040 36601 21098 36613
rect 21298 36789 21356 36801
rect 21298 36613 21310 36789
rect 21344 36613 21356 36789
rect 21298 36601 21356 36613
rect 21556 36789 21614 36801
rect 21556 36613 21568 36789
rect 21602 36613 21614 36789
rect 21556 36601 21614 36613
rect 21814 36789 21872 36801
rect 21814 36613 21826 36789
rect 21860 36613 21872 36789
rect 21814 36601 21872 36613
rect 22072 36789 22130 36801
rect 22072 36613 22084 36789
rect 22118 36613 22130 36789
rect 22072 36601 22130 36613
rect 22330 36789 22388 36801
rect 22330 36613 22342 36789
rect 22376 36613 22388 36789
rect 22330 36601 22388 36613
rect 22588 36789 22646 36801
rect 22588 36613 22600 36789
rect 22634 36613 22646 36789
rect 22588 36601 22646 36613
rect 22846 36789 22904 36801
rect 22846 36613 22858 36789
rect 22892 36613 22904 36789
rect 22846 36601 22904 36613
rect 23104 36789 23162 36801
rect 23104 36613 23116 36789
rect 23150 36613 23162 36789
rect 23104 36601 23162 36613
rect 23362 36789 23420 36801
rect 23362 36613 23374 36789
rect 23408 36613 23420 36789
rect 23362 36601 23420 36613
rect 20266 36353 20324 36365
rect 20266 36293 20278 36353
rect 20312 36293 20324 36353
rect 20266 36281 20324 36293
rect 20524 36353 20582 36365
rect 20524 36293 20536 36353
rect 20570 36293 20582 36353
rect 20524 36281 20582 36293
rect 20782 36353 20840 36365
rect 20782 36293 20794 36353
rect 20828 36293 20840 36353
rect 20782 36281 20840 36293
rect 21040 36353 21098 36365
rect 21040 36293 21052 36353
rect 21086 36293 21098 36353
rect 21040 36281 21098 36293
rect 21298 36353 21356 36365
rect 21298 36293 21310 36353
rect 21344 36293 21356 36353
rect 21298 36281 21356 36293
rect 21556 36353 21614 36365
rect 21556 36293 21568 36353
rect 21602 36293 21614 36353
rect 21556 36281 21614 36293
rect 21814 36353 21872 36365
rect 21814 36293 21826 36353
rect 21860 36293 21872 36353
rect 21814 36281 21872 36293
rect 22072 36353 22130 36365
rect 22072 36293 22084 36353
rect 22118 36293 22130 36353
rect 22072 36281 22130 36293
rect 22330 36353 22388 36365
rect 22330 36293 22342 36353
rect 22376 36293 22388 36353
rect 22330 36281 22388 36293
rect 22588 36353 22646 36365
rect 22588 36293 22600 36353
rect 22634 36293 22646 36353
rect 22588 36281 22646 36293
rect 22846 36353 22904 36365
rect 22846 36293 22858 36353
rect 22892 36293 22904 36353
rect 22846 36281 22904 36293
rect 23104 36353 23162 36365
rect 23104 36293 23116 36353
rect 23150 36293 23162 36353
rect 23104 36281 23162 36293
rect 23362 36353 23420 36365
rect 23362 36293 23374 36353
rect 23408 36293 23420 36353
rect 23362 36281 23420 36293
rect 12614 34999 12666 35083
rect 12614 34965 12622 34999
rect 12656 34965 12666 34999
rect 12614 34953 12666 34965
rect 12696 35067 12750 35083
rect 12696 35033 12706 35067
rect 12740 35033 12750 35067
rect 12696 34999 12750 35033
rect 12696 34965 12706 34999
rect 12740 34965 12750 34999
rect 12696 34953 12750 34965
rect 12780 34999 12834 35083
rect 12780 34965 12790 34999
rect 12824 34965 12834 34999
rect 12780 34953 12834 34965
rect 12864 35067 12918 35083
rect 12864 35033 12874 35067
rect 12908 35033 12918 35067
rect 12864 34999 12918 35033
rect 12864 34965 12874 34999
rect 12908 34965 12918 34999
rect 12864 34953 12918 34965
rect 12948 34999 13002 35083
rect 12948 34965 12958 34999
rect 12992 34965 13002 34999
rect 12948 34953 13002 34965
rect 13032 35067 13086 35083
rect 13032 35033 13042 35067
rect 13076 35033 13086 35067
rect 13032 34999 13086 35033
rect 13032 34965 13042 34999
rect 13076 34965 13086 34999
rect 13032 34953 13086 34965
rect 13116 34999 13170 35083
rect 13116 34965 13126 34999
rect 13160 34965 13170 34999
rect 13116 34953 13170 34965
rect 13200 35067 13254 35083
rect 13200 35033 13210 35067
rect 13244 35033 13254 35067
rect 13200 34999 13254 35033
rect 13200 34965 13210 34999
rect 13244 34965 13254 34999
rect 13200 34953 13254 34965
rect 13284 34999 13336 35083
rect 13284 34965 13294 34999
rect 13328 34965 13336 34999
rect 13284 34953 13336 34965
rect 25649 37921 25707 37933
rect 25649 37745 25661 37921
rect 25695 37745 25707 37921
rect 25649 37733 25707 37745
rect 25907 37921 25965 37933
rect 25907 37745 25919 37921
rect 25953 37745 25965 37921
rect 25907 37733 25965 37745
rect 26165 37921 26223 37933
rect 26165 37745 26177 37921
rect 26211 37745 26223 37921
rect 26165 37733 26223 37745
rect 25649 36461 25707 36473
rect 25649 36285 25661 36461
rect 25695 36285 25707 36461
rect 25649 36273 25707 36285
rect 25907 36461 25965 36473
rect 25907 36285 25919 36461
rect 25953 36285 25965 36461
rect 25907 36273 25965 36285
rect 26165 36461 26223 36473
rect 26165 36285 26177 36461
rect 26211 36285 26223 36461
rect 26165 36273 26223 36285
rect 25402 35117 25454 35201
rect 25402 35083 25410 35117
rect 25444 35083 25454 35117
rect 25402 35071 25454 35083
rect 25484 35185 25538 35201
rect 25484 35151 25494 35185
rect 25528 35151 25538 35185
rect 25484 35117 25538 35151
rect 25484 35083 25494 35117
rect 25528 35083 25538 35117
rect 25484 35071 25538 35083
rect 25568 35117 25622 35201
rect 25568 35083 25578 35117
rect 25612 35083 25622 35117
rect 25568 35071 25622 35083
rect 25652 35185 25706 35201
rect 25652 35151 25662 35185
rect 25696 35151 25706 35185
rect 25652 35117 25706 35151
rect 25652 35083 25662 35117
rect 25696 35083 25706 35117
rect 25652 35071 25706 35083
rect 25736 35117 25790 35201
rect 25736 35083 25746 35117
rect 25780 35083 25790 35117
rect 25736 35071 25790 35083
rect 25820 35185 25874 35201
rect 25820 35151 25830 35185
rect 25864 35151 25874 35185
rect 25820 35117 25874 35151
rect 25820 35083 25830 35117
rect 25864 35083 25874 35117
rect 25820 35071 25874 35083
rect 25904 35117 25958 35201
rect 25904 35083 25914 35117
rect 25948 35083 25958 35117
rect 25904 35071 25958 35083
rect 25988 35185 26042 35201
rect 25988 35151 25998 35185
rect 26032 35151 26042 35185
rect 25988 35117 26042 35151
rect 25988 35083 25998 35117
rect 26032 35083 26042 35117
rect 25988 35071 26042 35083
rect 26072 35117 26124 35201
rect 26072 35083 26082 35117
rect 26116 35083 26124 35117
rect 26072 35071 26124 35083
rect 7498 30745 7556 30757
rect 7498 30569 7510 30745
rect 7544 30569 7556 30745
rect 7498 30557 7556 30569
rect 7756 30745 7814 30757
rect 7756 30569 7768 30745
rect 7802 30569 7814 30745
rect 7756 30557 7814 30569
rect 8014 30745 8072 30757
rect 8014 30569 8026 30745
rect 8060 30569 8072 30745
rect 8014 30557 8072 30569
rect 8272 30745 8330 30757
rect 8272 30569 8284 30745
rect 8318 30569 8330 30745
rect 8272 30557 8330 30569
rect 8530 30745 8588 30757
rect 8530 30569 8542 30745
rect 8576 30569 8588 30745
rect 8530 30557 8588 30569
rect 8788 30745 8846 30757
rect 8788 30569 8800 30745
rect 8834 30569 8846 30745
rect 8788 30557 8846 30569
rect 9046 30745 9104 30757
rect 9046 30569 9058 30745
rect 9092 30569 9104 30745
rect 9046 30557 9104 30569
rect 9304 30745 9362 30757
rect 9304 30569 9316 30745
rect 9350 30569 9362 30745
rect 9304 30557 9362 30569
rect 9562 30745 9620 30757
rect 9562 30569 9574 30745
rect 9608 30569 9620 30745
rect 9562 30557 9620 30569
rect 9820 30745 9878 30757
rect 9820 30569 9832 30745
rect 9866 30569 9878 30745
rect 9820 30557 9878 30569
rect 10078 30745 10136 30757
rect 10078 30569 10090 30745
rect 10124 30569 10136 30745
rect 10078 30557 10136 30569
rect 10336 30745 10394 30757
rect 10336 30569 10348 30745
rect 10382 30569 10394 30745
rect 10336 30557 10394 30569
rect 10594 30745 10652 30757
rect 10594 30569 10606 30745
rect 10640 30569 10652 30745
rect 10594 30557 10652 30569
rect 7498 30309 7556 30321
rect 7498 30249 7510 30309
rect 7544 30249 7556 30309
rect 7498 30237 7556 30249
rect 7756 30309 7814 30321
rect 7756 30249 7768 30309
rect 7802 30249 7814 30309
rect 7756 30237 7814 30249
rect 8014 30309 8072 30321
rect 8014 30249 8026 30309
rect 8060 30249 8072 30309
rect 8014 30237 8072 30249
rect 8272 30309 8330 30321
rect 8272 30249 8284 30309
rect 8318 30249 8330 30309
rect 8272 30237 8330 30249
rect 8530 30309 8588 30321
rect 8530 30249 8542 30309
rect 8576 30249 8588 30309
rect 8530 30237 8588 30249
rect 8788 30309 8846 30321
rect 8788 30249 8800 30309
rect 8834 30249 8846 30309
rect 8788 30237 8846 30249
rect 9046 30309 9104 30321
rect 9046 30249 9058 30309
rect 9092 30249 9104 30309
rect 9046 30237 9104 30249
rect 9304 30309 9362 30321
rect 9304 30249 9316 30309
rect 9350 30249 9362 30309
rect 9304 30237 9362 30249
rect 9562 30309 9620 30321
rect 9562 30249 9574 30309
rect 9608 30249 9620 30309
rect 9562 30237 9620 30249
rect 9820 30309 9878 30321
rect 9820 30249 9832 30309
rect 9866 30249 9878 30309
rect 9820 30237 9878 30249
rect 10078 30309 10136 30321
rect 10078 30249 10090 30309
rect 10124 30249 10136 30309
rect 10078 30237 10136 30249
rect 10336 30309 10394 30321
rect 10336 30249 10348 30309
rect 10382 30249 10394 30309
rect 10336 30237 10394 30249
rect 10594 30309 10652 30321
rect 10594 30249 10606 30309
rect 10640 30249 10652 30309
rect 10594 30237 10652 30249
rect 12881 31877 12939 31889
rect 12881 31701 12893 31877
rect 12927 31701 12939 31877
rect 12881 31689 12939 31701
rect 13139 31877 13197 31889
rect 13139 31701 13151 31877
rect 13185 31701 13197 31877
rect 13139 31689 13197 31701
rect 13397 31877 13455 31889
rect 13397 31701 13409 31877
rect 13443 31701 13455 31877
rect 13397 31689 13455 31701
rect 12881 30417 12939 30429
rect 12881 30241 12893 30417
rect 12927 30241 12939 30417
rect 12881 30229 12939 30241
rect 13139 30417 13197 30429
rect 13139 30241 13151 30417
rect 13185 30241 13197 30417
rect 13139 30229 13197 30241
rect 13397 30417 13455 30429
rect 13397 30241 13409 30417
rect 13443 30241 13455 30417
rect 13397 30229 13455 30241
rect 20230 30669 20288 30681
rect 20230 30493 20242 30669
rect 20276 30493 20288 30669
rect 20230 30481 20288 30493
rect 20488 30669 20546 30681
rect 20488 30493 20500 30669
rect 20534 30493 20546 30669
rect 20488 30481 20546 30493
rect 20746 30669 20804 30681
rect 20746 30493 20758 30669
rect 20792 30493 20804 30669
rect 20746 30481 20804 30493
rect 21004 30669 21062 30681
rect 21004 30493 21016 30669
rect 21050 30493 21062 30669
rect 21004 30481 21062 30493
rect 21262 30669 21320 30681
rect 21262 30493 21274 30669
rect 21308 30493 21320 30669
rect 21262 30481 21320 30493
rect 21520 30669 21578 30681
rect 21520 30493 21532 30669
rect 21566 30493 21578 30669
rect 21520 30481 21578 30493
rect 21778 30669 21836 30681
rect 21778 30493 21790 30669
rect 21824 30493 21836 30669
rect 21778 30481 21836 30493
rect 22036 30669 22094 30681
rect 22036 30493 22048 30669
rect 22082 30493 22094 30669
rect 22036 30481 22094 30493
rect 22294 30669 22352 30681
rect 22294 30493 22306 30669
rect 22340 30493 22352 30669
rect 22294 30481 22352 30493
rect 22552 30669 22610 30681
rect 22552 30493 22564 30669
rect 22598 30493 22610 30669
rect 22552 30481 22610 30493
rect 22810 30669 22868 30681
rect 22810 30493 22822 30669
rect 22856 30493 22868 30669
rect 22810 30481 22868 30493
rect 23068 30669 23126 30681
rect 23068 30493 23080 30669
rect 23114 30493 23126 30669
rect 23068 30481 23126 30493
rect 23326 30669 23384 30681
rect 23326 30493 23338 30669
rect 23372 30493 23384 30669
rect 23326 30481 23384 30493
rect 20230 30233 20288 30245
rect 20230 30173 20242 30233
rect 20276 30173 20288 30233
rect 20230 30161 20288 30173
rect 20488 30233 20546 30245
rect 20488 30173 20500 30233
rect 20534 30173 20546 30233
rect 20488 30161 20546 30173
rect 20746 30233 20804 30245
rect 20746 30173 20758 30233
rect 20792 30173 20804 30233
rect 20746 30161 20804 30173
rect 21004 30233 21062 30245
rect 21004 30173 21016 30233
rect 21050 30173 21062 30233
rect 21004 30161 21062 30173
rect 21262 30233 21320 30245
rect 21262 30173 21274 30233
rect 21308 30173 21320 30233
rect 21262 30161 21320 30173
rect 21520 30233 21578 30245
rect 21520 30173 21532 30233
rect 21566 30173 21578 30233
rect 21520 30161 21578 30173
rect 21778 30233 21836 30245
rect 21778 30173 21790 30233
rect 21824 30173 21836 30233
rect 21778 30161 21836 30173
rect 22036 30233 22094 30245
rect 22036 30173 22048 30233
rect 22082 30173 22094 30233
rect 22036 30161 22094 30173
rect 22294 30233 22352 30245
rect 22294 30173 22306 30233
rect 22340 30173 22352 30233
rect 22294 30161 22352 30173
rect 22552 30233 22610 30245
rect 22552 30173 22564 30233
rect 22598 30173 22610 30233
rect 22552 30161 22610 30173
rect 22810 30233 22868 30245
rect 22810 30173 22822 30233
rect 22856 30173 22868 30233
rect 22810 30161 22868 30173
rect 23068 30233 23126 30245
rect 23068 30173 23080 30233
rect 23114 30173 23126 30233
rect 23068 30161 23126 30173
rect 23326 30233 23384 30245
rect 23326 30173 23338 30233
rect 23372 30173 23384 30233
rect 23326 30161 23384 30173
rect 12634 29073 12686 29157
rect 12634 29039 12642 29073
rect 12676 29039 12686 29073
rect 12634 29027 12686 29039
rect 12716 29141 12770 29157
rect 12716 29107 12726 29141
rect 12760 29107 12770 29141
rect 12716 29073 12770 29107
rect 12716 29039 12726 29073
rect 12760 29039 12770 29073
rect 12716 29027 12770 29039
rect 12800 29073 12854 29157
rect 12800 29039 12810 29073
rect 12844 29039 12854 29073
rect 12800 29027 12854 29039
rect 12884 29141 12938 29157
rect 12884 29107 12894 29141
rect 12928 29107 12938 29141
rect 12884 29073 12938 29107
rect 12884 29039 12894 29073
rect 12928 29039 12938 29073
rect 12884 29027 12938 29039
rect 12968 29073 13022 29157
rect 12968 29039 12978 29073
rect 13012 29039 13022 29073
rect 12968 29027 13022 29039
rect 13052 29141 13106 29157
rect 13052 29107 13062 29141
rect 13096 29107 13106 29141
rect 13052 29073 13106 29107
rect 13052 29039 13062 29073
rect 13096 29039 13106 29073
rect 13052 29027 13106 29039
rect 13136 29073 13190 29157
rect 13136 29039 13146 29073
rect 13180 29039 13190 29073
rect 13136 29027 13190 29039
rect 13220 29141 13274 29157
rect 13220 29107 13230 29141
rect 13264 29107 13274 29141
rect 13220 29073 13274 29107
rect 13220 29039 13230 29073
rect 13264 29039 13274 29073
rect 13220 29027 13274 29039
rect 13304 29073 13356 29157
rect 13304 29039 13314 29073
rect 13348 29039 13356 29073
rect 13304 29027 13356 29039
rect 25613 31801 25671 31813
rect 25613 31625 25625 31801
rect 25659 31625 25671 31801
rect 25613 31613 25671 31625
rect 25871 31801 25929 31813
rect 25871 31625 25883 31801
rect 25917 31625 25929 31801
rect 25871 31613 25929 31625
rect 26129 31801 26187 31813
rect 26129 31625 26141 31801
rect 26175 31625 26187 31801
rect 26129 31613 26187 31625
rect 25613 30341 25671 30353
rect 25613 30165 25625 30341
rect 25659 30165 25671 30341
rect 25613 30153 25671 30165
rect 25871 30341 25929 30353
rect 25871 30165 25883 30341
rect 25917 30165 25929 30341
rect 25871 30153 25929 30165
rect 26129 30341 26187 30353
rect 26129 30165 26141 30341
rect 26175 30165 26187 30341
rect 26129 30153 26187 30165
rect 25366 28997 25418 29081
rect 25366 28963 25374 28997
rect 25408 28963 25418 28997
rect 25366 28951 25418 28963
rect 25448 29065 25502 29081
rect 25448 29031 25458 29065
rect 25492 29031 25502 29065
rect 25448 28997 25502 29031
rect 25448 28963 25458 28997
rect 25492 28963 25502 28997
rect 25448 28951 25502 28963
rect 25532 28997 25586 29081
rect 25532 28963 25542 28997
rect 25576 28963 25586 28997
rect 25532 28951 25586 28963
rect 25616 29065 25670 29081
rect 25616 29031 25626 29065
rect 25660 29031 25670 29065
rect 25616 28997 25670 29031
rect 25616 28963 25626 28997
rect 25660 28963 25670 28997
rect 25616 28951 25670 28963
rect 25700 28997 25754 29081
rect 25700 28963 25710 28997
rect 25744 28963 25754 28997
rect 25700 28951 25754 28963
rect 25784 29065 25838 29081
rect 25784 29031 25794 29065
rect 25828 29031 25838 29065
rect 25784 28997 25838 29031
rect 25784 28963 25794 28997
rect 25828 28963 25838 28997
rect 25784 28951 25838 28963
rect 25868 28997 25922 29081
rect 25868 28963 25878 28997
rect 25912 28963 25922 28997
rect 25868 28951 25922 28963
rect 25952 29065 26006 29081
rect 25952 29031 25962 29065
rect 25996 29031 26006 29065
rect 25952 28997 26006 29031
rect 25952 28963 25962 28997
rect 25996 28963 26006 28997
rect 25952 28951 26006 28963
rect 26036 28997 26088 29081
rect 26036 28963 26046 28997
rect 26080 28963 26088 28997
rect 26036 28951 26088 28963
rect 7618 24041 7676 24053
rect 7618 23865 7630 24041
rect 7664 23865 7676 24041
rect 7618 23853 7676 23865
rect 7876 24041 7934 24053
rect 7876 23865 7888 24041
rect 7922 23865 7934 24041
rect 7876 23853 7934 23865
rect 8134 24041 8192 24053
rect 8134 23865 8146 24041
rect 8180 23865 8192 24041
rect 8134 23853 8192 23865
rect 8392 24041 8450 24053
rect 8392 23865 8404 24041
rect 8438 23865 8450 24041
rect 8392 23853 8450 23865
rect 8650 24041 8708 24053
rect 8650 23865 8662 24041
rect 8696 23865 8708 24041
rect 8650 23853 8708 23865
rect 8908 24041 8966 24053
rect 8908 23865 8920 24041
rect 8954 23865 8966 24041
rect 8908 23853 8966 23865
rect 9166 24041 9224 24053
rect 9166 23865 9178 24041
rect 9212 23865 9224 24041
rect 9166 23853 9224 23865
rect 9424 24041 9482 24053
rect 9424 23865 9436 24041
rect 9470 23865 9482 24041
rect 9424 23853 9482 23865
rect 9682 24041 9740 24053
rect 9682 23865 9694 24041
rect 9728 23865 9740 24041
rect 9682 23853 9740 23865
rect 9940 24041 9998 24053
rect 9940 23865 9952 24041
rect 9986 23865 9998 24041
rect 9940 23853 9998 23865
rect 10198 24041 10256 24053
rect 10198 23865 10210 24041
rect 10244 23865 10256 24041
rect 10198 23853 10256 23865
rect 10456 24041 10514 24053
rect 10456 23865 10468 24041
rect 10502 23865 10514 24041
rect 10456 23853 10514 23865
rect 10714 24041 10772 24053
rect 10714 23865 10726 24041
rect 10760 23865 10772 24041
rect 10714 23853 10772 23865
rect 7618 23605 7676 23617
rect 7618 23545 7630 23605
rect 7664 23545 7676 23605
rect 7618 23533 7676 23545
rect 7876 23605 7934 23617
rect 7876 23545 7888 23605
rect 7922 23545 7934 23605
rect 7876 23533 7934 23545
rect 8134 23605 8192 23617
rect 8134 23545 8146 23605
rect 8180 23545 8192 23605
rect 8134 23533 8192 23545
rect 8392 23605 8450 23617
rect 8392 23545 8404 23605
rect 8438 23545 8450 23605
rect 8392 23533 8450 23545
rect 8650 23605 8708 23617
rect 8650 23545 8662 23605
rect 8696 23545 8708 23605
rect 8650 23533 8708 23545
rect 8908 23605 8966 23617
rect 8908 23545 8920 23605
rect 8954 23545 8966 23605
rect 8908 23533 8966 23545
rect 9166 23605 9224 23617
rect 9166 23545 9178 23605
rect 9212 23545 9224 23605
rect 9166 23533 9224 23545
rect 9424 23605 9482 23617
rect 9424 23545 9436 23605
rect 9470 23545 9482 23605
rect 9424 23533 9482 23545
rect 9682 23605 9740 23617
rect 9682 23545 9694 23605
rect 9728 23545 9740 23605
rect 9682 23533 9740 23545
rect 9940 23605 9998 23617
rect 9940 23545 9952 23605
rect 9986 23545 9998 23605
rect 9940 23533 9998 23545
rect 10198 23605 10256 23617
rect 10198 23545 10210 23605
rect 10244 23545 10256 23605
rect 10198 23533 10256 23545
rect 10456 23605 10514 23617
rect 10456 23545 10468 23605
rect 10502 23545 10514 23605
rect 10456 23533 10514 23545
rect 10714 23605 10772 23617
rect 10714 23545 10726 23605
rect 10760 23545 10772 23605
rect 10714 23533 10772 23545
rect 13001 25173 13059 25185
rect 13001 24997 13013 25173
rect 13047 24997 13059 25173
rect 13001 24985 13059 24997
rect 13259 25173 13317 25185
rect 13259 24997 13271 25173
rect 13305 24997 13317 25173
rect 13259 24985 13317 24997
rect 13517 25173 13575 25185
rect 13517 24997 13529 25173
rect 13563 24997 13575 25173
rect 13517 24985 13575 24997
rect 13001 23713 13059 23725
rect 13001 23537 13013 23713
rect 13047 23537 13059 23713
rect 13001 23525 13059 23537
rect 13259 23713 13317 23725
rect 13259 23537 13271 23713
rect 13305 23537 13317 23713
rect 13259 23525 13317 23537
rect 13517 23713 13575 23725
rect 13517 23537 13529 23713
rect 13563 23537 13575 23713
rect 13517 23525 13575 23537
rect 20326 23911 20384 23923
rect 20326 23735 20338 23911
rect 20372 23735 20384 23911
rect 20326 23723 20384 23735
rect 20584 23911 20642 23923
rect 20584 23735 20596 23911
rect 20630 23735 20642 23911
rect 20584 23723 20642 23735
rect 20842 23911 20900 23923
rect 20842 23735 20854 23911
rect 20888 23735 20900 23911
rect 20842 23723 20900 23735
rect 21100 23911 21158 23923
rect 21100 23735 21112 23911
rect 21146 23735 21158 23911
rect 21100 23723 21158 23735
rect 21358 23911 21416 23923
rect 21358 23735 21370 23911
rect 21404 23735 21416 23911
rect 21358 23723 21416 23735
rect 21616 23911 21674 23923
rect 21616 23735 21628 23911
rect 21662 23735 21674 23911
rect 21616 23723 21674 23735
rect 21874 23911 21932 23923
rect 21874 23735 21886 23911
rect 21920 23735 21932 23911
rect 21874 23723 21932 23735
rect 22132 23911 22190 23923
rect 22132 23735 22144 23911
rect 22178 23735 22190 23911
rect 22132 23723 22190 23735
rect 22390 23911 22448 23923
rect 22390 23735 22402 23911
rect 22436 23735 22448 23911
rect 22390 23723 22448 23735
rect 22648 23911 22706 23923
rect 22648 23735 22660 23911
rect 22694 23735 22706 23911
rect 22648 23723 22706 23735
rect 22906 23911 22964 23923
rect 22906 23735 22918 23911
rect 22952 23735 22964 23911
rect 22906 23723 22964 23735
rect 23164 23911 23222 23923
rect 23164 23735 23176 23911
rect 23210 23735 23222 23911
rect 23164 23723 23222 23735
rect 23422 23911 23480 23923
rect 23422 23735 23434 23911
rect 23468 23735 23480 23911
rect 23422 23723 23480 23735
rect 20326 23475 20384 23487
rect 20326 23415 20338 23475
rect 20372 23415 20384 23475
rect 20326 23403 20384 23415
rect 20584 23475 20642 23487
rect 20584 23415 20596 23475
rect 20630 23415 20642 23475
rect 20584 23403 20642 23415
rect 20842 23475 20900 23487
rect 20842 23415 20854 23475
rect 20888 23415 20900 23475
rect 20842 23403 20900 23415
rect 21100 23475 21158 23487
rect 21100 23415 21112 23475
rect 21146 23415 21158 23475
rect 21100 23403 21158 23415
rect 21358 23475 21416 23487
rect 21358 23415 21370 23475
rect 21404 23415 21416 23475
rect 21358 23403 21416 23415
rect 21616 23475 21674 23487
rect 21616 23415 21628 23475
rect 21662 23415 21674 23475
rect 21616 23403 21674 23415
rect 21874 23475 21932 23487
rect 21874 23415 21886 23475
rect 21920 23415 21932 23475
rect 21874 23403 21932 23415
rect 22132 23475 22190 23487
rect 22132 23415 22144 23475
rect 22178 23415 22190 23475
rect 22132 23403 22190 23415
rect 22390 23475 22448 23487
rect 22390 23415 22402 23475
rect 22436 23415 22448 23475
rect 22390 23403 22448 23415
rect 22648 23475 22706 23487
rect 22648 23415 22660 23475
rect 22694 23415 22706 23475
rect 22648 23403 22706 23415
rect 22906 23475 22964 23487
rect 22906 23415 22918 23475
rect 22952 23415 22964 23475
rect 22906 23403 22964 23415
rect 23164 23475 23222 23487
rect 23164 23415 23176 23475
rect 23210 23415 23222 23475
rect 23164 23403 23222 23415
rect 23422 23475 23480 23487
rect 23422 23415 23434 23475
rect 23468 23415 23480 23475
rect 23422 23403 23480 23415
rect 12754 22369 12806 22453
rect 12754 22335 12762 22369
rect 12796 22335 12806 22369
rect 12754 22323 12806 22335
rect 12836 22437 12890 22453
rect 12836 22403 12846 22437
rect 12880 22403 12890 22437
rect 12836 22369 12890 22403
rect 12836 22335 12846 22369
rect 12880 22335 12890 22369
rect 12836 22323 12890 22335
rect 12920 22369 12974 22453
rect 12920 22335 12930 22369
rect 12964 22335 12974 22369
rect 12920 22323 12974 22335
rect 13004 22437 13058 22453
rect 13004 22403 13014 22437
rect 13048 22403 13058 22437
rect 13004 22369 13058 22403
rect 13004 22335 13014 22369
rect 13048 22335 13058 22369
rect 13004 22323 13058 22335
rect 13088 22369 13142 22453
rect 13088 22335 13098 22369
rect 13132 22335 13142 22369
rect 13088 22323 13142 22335
rect 13172 22437 13226 22453
rect 13172 22403 13182 22437
rect 13216 22403 13226 22437
rect 13172 22369 13226 22403
rect 13172 22335 13182 22369
rect 13216 22335 13226 22369
rect 13172 22323 13226 22335
rect 13256 22369 13310 22453
rect 13256 22335 13266 22369
rect 13300 22335 13310 22369
rect 13256 22323 13310 22335
rect 13340 22437 13394 22453
rect 13340 22403 13350 22437
rect 13384 22403 13394 22437
rect 13340 22369 13394 22403
rect 13340 22335 13350 22369
rect 13384 22335 13394 22369
rect 13340 22323 13394 22335
rect 13424 22369 13476 22453
rect 13424 22335 13434 22369
rect 13468 22335 13476 22369
rect 13424 22323 13476 22335
rect 25709 25043 25767 25055
rect 25709 24867 25721 25043
rect 25755 24867 25767 25043
rect 25709 24855 25767 24867
rect 25967 25043 26025 25055
rect 25967 24867 25979 25043
rect 26013 24867 26025 25043
rect 25967 24855 26025 24867
rect 26225 25043 26283 25055
rect 26225 24867 26237 25043
rect 26271 24867 26283 25043
rect 26225 24855 26283 24867
rect 25709 23583 25767 23595
rect 25709 23407 25721 23583
rect 25755 23407 25767 23583
rect 25709 23395 25767 23407
rect 25967 23583 26025 23595
rect 25967 23407 25979 23583
rect 26013 23407 26025 23583
rect 25967 23395 26025 23407
rect 26225 23583 26283 23595
rect 26225 23407 26237 23583
rect 26271 23407 26283 23583
rect 26225 23395 26283 23407
rect 25462 22239 25514 22323
rect 25462 22205 25470 22239
rect 25504 22205 25514 22239
rect 25462 22193 25514 22205
rect 25544 22307 25598 22323
rect 25544 22273 25554 22307
rect 25588 22273 25598 22307
rect 25544 22239 25598 22273
rect 25544 22205 25554 22239
rect 25588 22205 25598 22239
rect 25544 22193 25598 22205
rect 25628 22239 25682 22323
rect 25628 22205 25638 22239
rect 25672 22205 25682 22239
rect 25628 22193 25682 22205
rect 25712 22307 25766 22323
rect 25712 22273 25722 22307
rect 25756 22273 25766 22307
rect 25712 22239 25766 22273
rect 25712 22205 25722 22239
rect 25756 22205 25766 22239
rect 25712 22193 25766 22205
rect 25796 22239 25850 22323
rect 25796 22205 25806 22239
rect 25840 22205 25850 22239
rect 25796 22193 25850 22205
rect 25880 22307 25934 22323
rect 25880 22273 25890 22307
rect 25924 22273 25934 22307
rect 25880 22239 25934 22273
rect 25880 22205 25890 22239
rect 25924 22205 25934 22239
rect 25880 22193 25934 22205
rect 25964 22239 26018 22323
rect 25964 22205 25974 22239
rect 26008 22205 26018 22239
rect 25964 22193 26018 22205
rect 26048 22307 26102 22323
rect 26048 22273 26058 22307
rect 26092 22273 26102 22307
rect 26048 22239 26102 22273
rect 26048 22205 26058 22239
rect 26092 22205 26102 22239
rect 26048 22193 26102 22205
rect 26132 22239 26184 22323
rect 26132 22205 26142 22239
rect 26176 22205 26184 22239
rect 26132 22193 26184 22205
rect 7494 16995 7552 17007
rect 7494 16819 7506 16995
rect 7540 16819 7552 16995
rect 7494 16807 7552 16819
rect 7752 16995 7810 17007
rect 7752 16819 7764 16995
rect 7798 16819 7810 16995
rect 7752 16807 7810 16819
rect 8010 16995 8068 17007
rect 8010 16819 8022 16995
rect 8056 16819 8068 16995
rect 8010 16807 8068 16819
rect 8268 16995 8326 17007
rect 8268 16819 8280 16995
rect 8314 16819 8326 16995
rect 8268 16807 8326 16819
rect 8526 16995 8584 17007
rect 8526 16819 8538 16995
rect 8572 16819 8584 16995
rect 8526 16807 8584 16819
rect 8784 16995 8842 17007
rect 8784 16819 8796 16995
rect 8830 16819 8842 16995
rect 8784 16807 8842 16819
rect 9042 16995 9100 17007
rect 9042 16819 9054 16995
rect 9088 16819 9100 16995
rect 9042 16807 9100 16819
rect 9300 16995 9358 17007
rect 9300 16819 9312 16995
rect 9346 16819 9358 16995
rect 9300 16807 9358 16819
rect 9558 16995 9616 17007
rect 9558 16819 9570 16995
rect 9604 16819 9616 16995
rect 9558 16807 9616 16819
rect 9816 16995 9874 17007
rect 9816 16819 9828 16995
rect 9862 16819 9874 16995
rect 9816 16807 9874 16819
rect 10074 16995 10132 17007
rect 10074 16819 10086 16995
rect 10120 16819 10132 16995
rect 10074 16807 10132 16819
rect 10332 16995 10390 17007
rect 10332 16819 10344 16995
rect 10378 16819 10390 16995
rect 10332 16807 10390 16819
rect 10590 16995 10648 17007
rect 10590 16819 10602 16995
rect 10636 16819 10648 16995
rect 10590 16807 10648 16819
rect 7494 16559 7552 16571
rect 7494 16499 7506 16559
rect 7540 16499 7552 16559
rect 7494 16487 7552 16499
rect 7752 16559 7810 16571
rect 7752 16499 7764 16559
rect 7798 16499 7810 16559
rect 7752 16487 7810 16499
rect 8010 16559 8068 16571
rect 8010 16499 8022 16559
rect 8056 16499 8068 16559
rect 8010 16487 8068 16499
rect 8268 16559 8326 16571
rect 8268 16499 8280 16559
rect 8314 16499 8326 16559
rect 8268 16487 8326 16499
rect 8526 16559 8584 16571
rect 8526 16499 8538 16559
rect 8572 16499 8584 16559
rect 8526 16487 8584 16499
rect 8784 16559 8842 16571
rect 8784 16499 8796 16559
rect 8830 16499 8842 16559
rect 8784 16487 8842 16499
rect 9042 16559 9100 16571
rect 9042 16499 9054 16559
rect 9088 16499 9100 16559
rect 9042 16487 9100 16499
rect 9300 16559 9358 16571
rect 9300 16499 9312 16559
rect 9346 16499 9358 16559
rect 9300 16487 9358 16499
rect 9558 16559 9616 16571
rect 9558 16499 9570 16559
rect 9604 16499 9616 16559
rect 9558 16487 9616 16499
rect 9816 16559 9874 16571
rect 9816 16499 9828 16559
rect 9862 16499 9874 16559
rect 9816 16487 9874 16499
rect 10074 16559 10132 16571
rect 10074 16499 10086 16559
rect 10120 16499 10132 16559
rect 10074 16487 10132 16499
rect 10332 16559 10390 16571
rect 10332 16499 10344 16559
rect 10378 16499 10390 16559
rect 10332 16487 10390 16499
rect 10590 16559 10648 16571
rect 10590 16499 10602 16559
rect 10636 16499 10648 16559
rect 10590 16487 10648 16499
rect 12877 18127 12935 18139
rect 12877 17951 12889 18127
rect 12923 17951 12935 18127
rect 12877 17939 12935 17951
rect 13135 18127 13193 18139
rect 13135 17951 13147 18127
rect 13181 17951 13193 18127
rect 13135 17939 13193 17951
rect 13393 18127 13451 18139
rect 13393 17951 13405 18127
rect 13439 17951 13451 18127
rect 13393 17939 13451 17951
rect 12877 16667 12935 16679
rect 12877 16491 12889 16667
rect 12923 16491 12935 16667
rect 12877 16479 12935 16491
rect 13135 16667 13193 16679
rect 13135 16491 13147 16667
rect 13181 16491 13193 16667
rect 13135 16479 13193 16491
rect 13393 16667 13451 16679
rect 13393 16491 13405 16667
rect 13439 16491 13451 16667
rect 13393 16479 13451 16491
rect 20676 16865 20734 16877
rect 20676 16689 20688 16865
rect 20722 16689 20734 16865
rect 20676 16677 20734 16689
rect 20934 16865 20992 16877
rect 20934 16689 20946 16865
rect 20980 16689 20992 16865
rect 20934 16677 20992 16689
rect 21192 16865 21250 16877
rect 21192 16689 21204 16865
rect 21238 16689 21250 16865
rect 21192 16677 21250 16689
rect 21450 16865 21508 16877
rect 21450 16689 21462 16865
rect 21496 16689 21508 16865
rect 21450 16677 21508 16689
rect 21708 16865 21766 16877
rect 21708 16689 21720 16865
rect 21754 16689 21766 16865
rect 21708 16677 21766 16689
rect 21966 16865 22024 16877
rect 21966 16689 21978 16865
rect 22012 16689 22024 16865
rect 21966 16677 22024 16689
rect 22224 16865 22282 16877
rect 22224 16689 22236 16865
rect 22270 16689 22282 16865
rect 22224 16677 22282 16689
rect 22482 16865 22540 16877
rect 22482 16689 22494 16865
rect 22528 16689 22540 16865
rect 22482 16677 22540 16689
rect 22740 16865 22798 16877
rect 22740 16689 22752 16865
rect 22786 16689 22798 16865
rect 22740 16677 22798 16689
rect 22998 16865 23056 16877
rect 22998 16689 23010 16865
rect 23044 16689 23056 16865
rect 22998 16677 23056 16689
rect 23256 16865 23314 16877
rect 23256 16689 23268 16865
rect 23302 16689 23314 16865
rect 23256 16677 23314 16689
rect 23514 16865 23572 16877
rect 23514 16689 23526 16865
rect 23560 16689 23572 16865
rect 23514 16677 23572 16689
rect 23772 16865 23830 16877
rect 23772 16689 23784 16865
rect 23818 16689 23830 16865
rect 23772 16677 23830 16689
rect 20676 16429 20734 16441
rect 20676 16369 20688 16429
rect 20722 16369 20734 16429
rect 20676 16357 20734 16369
rect 20934 16429 20992 16441
rect 20934 16369 20946 16429
rect 20980 16369 20992 16429
rect 20934 16357 20992 16369
rect 21192 16429 21250 16441
rect 21192 16369 21204 16429
rect 21238 16369 21250 16429
rect 21192 16357 21250 16369
rect 21450 16429 21508 16441
rect 21450 16369 21462 16429
rect 21496 16369 21508 16429
rect 21450 16357 21508 16369
rect 21708 16429 21766 16441
rect 21708 16369 21720 16429
rect 21754 16369 21766 16429
rect 21708 16357 21766 16369
rect 21966 16429 22024 16441
rect 21966 16369 21978 16429
rect 22012 16369 22024 16429
rect 21966 16357 22024 16369
rect 22224 16429 22282 16441
rect 22224 16369 22236 16429
rect 22270 16369 22282 16429
rect 22224 16357 22282 16369
rect 22482 16429 22540 16441
rect 22482 16369 22494 16429
rect 22528 16369 22540 16429
rect 22482 16357 22540 16369
rect 22740 16429 22798 16441
rect 22740 16369 22752 16429
rect 22786 16369 22798 16429
rect 22740 16357 22798 16369
rect 22998 16429 23056 16441
rect 22998 16369 23010 16429
rect 23044 16369 23056 16429
rect 22998 16357 23056 16369
rect 23256 16429 23314 16441
rect 23256 16369 23268 16429
rect 23302 16369 23314 16429
rect 23256 16357 23314 16369
rect 23514 16429 23572 16441
rect 23514 16369 23526 16429
rect 23560 16369 23572 16429
rect 23514 16357 23572 16369
rect 23772 16429 23830 16441
rect 23772 16369 23784 16429
rect 23818 16369 23830 16429
rect 23772 16357 23830 16369
rect 12630 15323 12682 15407
rect 12630 15289 12638 15323
rect 12672 15289 12682 15323
rect 12630 15277 12682 15289
rect 12712 15391 12766 15407
rect 12712 15357 12722 15391
rect 12756 15357 12766 15391
rect 12712 15323 12766 15357
rect 12712 15289 12722 15323
rect 12756 15289 12766 15323
rect 12712 15277 12766 15289
rect 12796 15323 12850 15407
rect 12796 15289 12806 15323
rect 12840 15289 12850 15323
rect 12796 15277 12850 15289
rect 12880 15391 12934 15407
rect 12880 15357 12890 15391
rect 12924 15357 12934 15391
rect 12880 15323 12934 15357
rect 12880 15289 12890 15323
rect 12924 15289 12934 15323
rect 12880 15277 12934 15289
rect 12964 15323 13018 15407
rect 12964 15289 12974 15323
rect 13008 15289 13018 15323
rect 12964 15277 13018 15289
rect 13048 15391 13102 15407
rect 13048 15357 13058 15391
rect 13092 15357 13102 15391
rect 13048 15323 13102 15357
rect 13048 15289 13058 15323
rect 13092 15289 13102 15323
rect 13048 15277 13102 15289
rect 13132 15323 13186 15407
rect 13132 15289 13142 15323
rect 13176 15289 13186 15323
rect 13132 15277 13186 15289
rect 13216 15391 13270 15407
rect 13216 15357 13226 15391
rect 13260 15357 13270 15391
rect 13216 15323 13270 15357
rect 13216 15289 13226 15323
rect 13260 15289 13270 15323
rect 13216 15277 13270 15289
rect 13300 15323 13352 15407
rect 13300 15289 13310 15323
rect 13344 15289 13352 15323
rect 13300 15277 13352 15289
rect 26059 17997 26117 18009
rect 26059 17821 26071 17997
rect 26105 17821 26117 17997
rect 26059 17809 26117 17821
rect 26317 17997 26375 18009
rect 26317 17821 26329 17997
rect 26363 17821 26375 17997
rect 26317 17809 26375 17821
rect 26575 17997 26633 18009
rect 26575 17821 26587 17997
rect 26621 17821 26633 17997
rect 26575 17809 26633 17821
rect 26059 16537 26117 16549
rect 26059 16361 26071 16537
rect 26105 16361 26117 16537
rect 26059 16349 26117 16361
rect 26317 16537 26375 16549
rect 26317 16361 26329 16537
rect 26363 16361 26375 16537
rect 26317 16349 26375 16361
rect 26575 16537 26633 16549
rect 26575 16361 26587 16537
rect 26621 16361 26633 16537
rect 26575 16349 26633 16361
rect 25812 15193 25864 15277
rect 25812 15159 25820 15193
rect 25854 15159 25864 15193
rect 25812 15147 25864 15159
rect 25894 15261 25948 15277
rect 25894 15227 25904 15261
rect 25938 15227 25948 15261
rect 25894 15193 25948 15227
rect 25894 15159 25904 15193
rect 25938 15159 25948 15193
rect 25894 15147 25948 15159
rect 25978 15193 26032 15277
rect 25978 15159 25988 15193
rect 26022 15159 26032 15193
rect 25978 15147 26032 15159
rect 26062 15261 26116 15277
rect 26062 15227 26072 15261
rect 26106 15227 26116 15261
rect 26062 15193 26116 15227
rect 26062 15159 26072 15193
rect 26106 15159 26116 15193
rect 26062 15147 26116 15159
rect 26146 15193 26200 15277
rect 26146 15159 26156 15193
rect 26190 15159 26200 15193
rect 26146 15147 26200 15159
rect 26230 15261 26284 15277
rect 26230 15227 26240 15261
rect 26274 15227 26284 15261
rect 26230 15193 26284 15227
rect 26230 15159 26240 15193
rect 26274 15159 26284 15193
rect 26230 15147 26284 15159
rect 26314 15193 26368 15277
rect 26314 15159 26324 15193
rect 26358 15159 26368 15193
rect 26314 15147 26368 15159
rect 26398 15261 26452 15277
rect 26398 15227 26408 15261
rect 26442 15227 26452 15261
rect 26398 15193 26452 15227
rect 26398 15159 26408 15193
rect 26442 15159 26452 15193
rect 26398 15147 26452 15159
rect 26482 15193 26534 15277
rect 26482 15159 26492 15193
rect 26526 15159 26534 15193
rect 26482 15147 26534 15159
<< pdiff >>
rect 12861 38299 12919 38311
rect 12861 38123 12873 38299
rect 12907 38123 12919 38299
rect 12861 38111 12919 38123
rect 13119 38299 13177 38311
rect 13119 38123 13131 38299
rect 13165 38123 13177 38299
rect 13119 38111 13177 38123
rect 13377 38299 13435 38311
rect 13377 38123 13389 38299
rect 13423 38123 13435 38299
rect 13377 38111 13435 38123
rect 25649 38417 25707 38429
rect 25649 38241 25661 38417
rect 25695 38241 25707 38417
rect 25649 38229 25707 38241
rect 25907 38417 25965 38429
rect 25907 38241 25919 38417
rect 25953 38241 25965 38417
rect 25907 38229 25965 38241
rect 26165 38417 26223 38429
rect 26165 38241 26177 38417
rect 26211 38241 26223 38417
rect 26165 38229 26223 38241
rect 7478 37098 7536 37110
rect 7478 36922 7490 37098
rect 7524 36922 7536 37098
rect 7478 36910 7536 36922
rect 7736 37098 7794 37110
rect 7736 36922 7748 37098
rect 7782 36922 7794 37098
rect 7736 36910 7794 36922
rect 7994 37098 8052 37110
rect 7994 36922 8006 37098
rect 8040 36922 8052 37098
rect 7994 36910 8052 36922
rect 8252 37098 8310 37110
rect 8252 36922 8264 37098
rect 8298 36922 8310 37098
rect 8252 36910 8310 36922
rect 8510 37098 8568 37110
rect 8510 36922 8522 37098
rect 8556 36922 8568 37098
rect 8510 36910 8568 36922
rect 8768 37098 8826 37110
rect 8768 36922 8780 37098
rect 8814 36922 8826 37098
rect 8768 36910 8826 36922
rect 9026 37098 9084 37110
rect 9026 36922 9038 37098
rect 9072 36922 9084 37098
rect 9026 36910 9084 36922
rect 9284 37098 9342 37110
rect 9284 36922 9296 37098
rect 9330 36922 9342 37098
rect 9284 36910 9342 36922
rect 9542 37098 9600 37110
rect 9542 36922 9554 37098
rect 9588 36922 9600 37098
rect 9542 36910 9600 36922
rect 9800 37098 9858 37110
rect 9800 36922 9812 37098
rect 9846 36922 9858 37098
rect 9800 36910 9858 36922
rect 10058 37098 10116 37110
rect 10058 36922 10070 37098
rect 10104 36922 10116 37098
rect 10058 36910 10116 36922
rect 10316 37098 10374 37110
rect 10316 36922 10328 37098
rect 10362 36922 10374 37098
rect 10316 36910 10374 36922
rect 10574 37098 10632 37110
rect 10574 36922 10586 37098
rect 10620 36922 10632 37098
rect 10574 36910 10632 36922
rect 12861 36839 12919 36851
rect 12861 36663 12873 36839
rect 12907 36663 12919 36839
rect 12861 36651 12919 36663
rect 13119 36839 13177 36851
rect 13119 36663 13131 36839
rect 13165 36663 13177 36839
rect 13119 36651 13177 36663
rect 13377 36839 13435 36851
rect 13377 36663 13389 36839
rect 13423 36663 13435 36839
rect 13377 36651 13435 36663
rect 20266 37216 20324 37228
rect 20266 37040 20278 37216
rect 20312 37040 20324 37216
rect 20266 37028 20324 37040
rect 20524 37216 20582 37228
rect 20524 37040 20536 37216
rect 20570 37040 20582 37216
rect 20524 37028 20582 37040
rect 20782 37216 20840 37228
rect 20782 37040 20794 37216
rect 20828 37040 20840 37216
rect 20782 37028 20840 37040
rect 21040 37216 21098 37228
rect 21040 37040 21052 37216
rect 21086 37040 21098 37216
rect 21040 37028 21098 37040
rect 21298 37216 21356 37228
rect 21298 37040 21310 37216
rect 21344 37040 21356 37216
rect 21298 37028 21356 37040
rect 21556 37216 21614 37228
rect 21556 37040 21568 37216
rect 21602 37040 21614 37216
rect 21556 37028 21614 37040
rect 21814 37216 21872 37228
rect 21814 37040 21826 37216
rect 21860 37040 21872 37216
rect 21814 37028 21872 37040
rect 22072 37216 22130 37228
rect 22072 37040 22084 37216
rect 22118 37040 22130 37216
rect 22072 37028 22130 37040
rect 22330 37216 22388 37228
rect 22330 37040 22342 37216
rect 22376 37040 22388 37216
rect 22330 37028 22388 37040
rect 22588 37216 22646 37228
rect 22588 37040 22600 37216
rect 22634 37040 22646 37216
rect 22588 37028 22646 37040
rect 22846 37216 22904 37228
rect 22846 37040 22858 37216
rect 22892 37040 22904 37216
rect 22846 37028 22904 37040
rect 23104 37216 23162 37228
rect 23104 37040 23116 37216
rect 23150 37040 23162 37216
rect 23104 37028 23162 37040
rect 23362 37216 23420 37228
rect 23362 37040 23374 37216
rect 23408 37040 23420 37216
rect 23362 37028 23420 37040
rect 12614 35391 12666 35403
rect 12614 35357 12622 35391
rect 12656 35357 12666 35391
rect 12614 35323 12666 35357
rect 12614 35289 12622 35323
rect 12656 35289 12666 35323
rect 12614 35203 12666 35289
rect 12696 35391 12750 35403
rect 12696 35357 12706 35391
rect 12740 35357 12750 35391
rect 12696 35323 12750 35357
rect 12696 35289 12706 35323
rect 12740 35289 12750 35323
rect 12696 35255 12750 35289
rect 12696 35221 12706 35255
rect 12740 35221 12750 35255
rect 12696 35203 12750 35221
rect 12780 35391 12834 35403
rect 12780 35357 12790 35391
rect 12824 35357 12834 35391
rect 12780 35323 12834 35357
rect 12780 35289 12790 35323
rect 12824 35289 12834 35323
rect 12780 35203 12834 35289
rect 12864 35391 12918 35403
rect 12864 35357 12874 35391
rect 12908 35357 12918 35391
rect 12864 35323 12918 35357
rect 12864 35289 12874 35323
rect 12908 35289 12918 35323
rect 12864 35255 12918 35289
rect 12864 35221 12874 35255
rect 12908 35221 12918 35255
rect 12864 35203 12918 35221
rect 12948 35391 13002 35403
rect 12948 35357 12958 35391
rect 12992 35357 13002 35391
rect 12948 35323 13002 35357
rect 12948 35289 12958 35323
rect 12992 35289 13002 35323
rect 12948 35203 13002 35289
rect 13032 35391 13086 35403
rect 13032 35357 13042 35391
rect 13076 35357 13086 35391
rect 13032 35323 13086 35357
rect 13032 35289 13042 35323
rect 13076 35289 13086 35323
rect 13032 35255 13086 35289
rect 13032 35221 13042 35255
rect 13076 35221 13086 35255
rect 13032 35203 13086 35221
rect 13116 35391 13170 35403
rect 13116 35357 13126 35391
rect 13160 35357 13170 35391
rect 13116 35323 13170 35357
rect 13116 35289 13126 35323
rect 13160 35289 13170 35323
rect 13116 35203 13170 35289
rect 13200 35391 13254 35403
rect 13200 35357 13210 35391
rect 13244 35357 13254 35391
rect 13200 35323 13254 35357
rect 13200 35289 13210 35323
rect 13244 35289 13254 35323
rect 13200 35255 13254 35289
rect 13200 35221 13210 35255
rect 13244 35221 13254 35255
rect 13200 35203 13254 35221
rect 13284 35391 13336 35403
rect 13284 35357 13294 35391
rect 13328 35357 13336 35391
rect 13284 35323 13336 35357
rect 13284 35289 13294 35323
rect 13328 35289 13336 35323
rect 13284 35203 13336 35289
rect 25649 36957 25707 36969
rect 25649 36781 25661 36957
rect 25695 36781 25707 36957
rect 25649 36769 25707 36781
rect 25907 36957 25965 36969
rect 25907 36781 25919 36957
rect 25953 36781 25965 36957
rect 25907 36769 25965 36781
rect 26165 36957 26223 36969
rect 26165 36781 26177 36957
rect 26211 36781 26223 36957
rect 26165 36769 26223 36781
rect 25402 35509 25454 35521
rect 25402 35475 25410 35509
rect 25444 35475 25454 35509
rect 25402 35441 25454 35475
rect 25402 35407 25410 35441
rect 25444 35407 25454 35441
rect 25402 35321 25454 35407
rect 25484 35509 25538 35521
rect 25484 35475 25494 35509
rect 25528 35475 25538 35509
rect 25484 35441 25538 35475
rect 25484 35407 25494 35441
rect 25528 35407 25538 35441
rect 25484 35373 25538 35407
rect 25484 35339 25494 35373
rect 25528 35339 25538 35373
rect 25484 35321 25538 35339
rect 25568 35509 25622 35521
rect 25568 35475 25578 35509
rect 25612 35475 25622 35509
rect 25568 35441 25622 35475
rect 25568 35407 25578 35441
rect 25612 35407 25622 35441
rect 25568 35321 25622 35407
rect 25652 35509 25706 35521
rect 25652 35475 25662 35509
rect 25696 35475 25706 35509
rect 25652 35441 25706 35475
rect 25652 35407 25662 35441
rect 25696 35407 25706 35441
rect 25652 35373 25706 35407
rect 25652 35339 25662 35373
rect 25696 35339 25706 35373
rect 25652 35321 25706 35339
rect 25736 35509 25790 35521
rect 25736 35475 25746 35509
rect 25780 35475 25790 35509
rect 25736 35441 25790 35475
rect 25736 35407 25746 35441
rect 25780 35407 25790 35441
rect 25736 35321 25790 35407
rect 25820 35509 25874 35521
rect 25820 35475 25830 35509
rect 25864 35475 25874 35509
rect 25820 35441 25874 35475
rect 25820 35407 25830 35441
rect 25864 35407 25874 35441
rect 25820 35373 25874 35407
rect 25820 35339 25830 35373
rect 25864 35339 25874 35373
rect 25820 35321 25874 35339
rect 25904 35509 25958 35521
rect 25904 35475 25914 35509
rect 25948 35475 25958 35509
rect 25904 35441 25958 35475
rect 25904 35407 25914 35441
rect 25948 35407 25958 35441
rect 25904 35321 25958 35407
rect 25988 35509 26042 35521
rect 25988 35475 25998 35509
rect 26032 35475 26042 35509
rect 25988 35441 26042 35475
rect 25988 35407 25998 35441
rect 26032 35407 26042 35441
rect 25988 35373 26042 35407
rect 25988 35339 25998 35373
rect 26032 35339 26042 35373
rect 25988 35321 26042 35339
rect 26072 35509 26124 35521
rect 26072 35475 26082 35509
rect 26116 35475 26124 35509
rect 26072 35441 26124 35475
rect 26072 35407 26082 35441
rect 26116 35407 26124 35441
rect 26072 35321 26124 35407
rect 12881 32373 12939 32385
rect 12881 32197 12893 32373
rect 12927 32197 12939 32373
rect 12881 32185 12939 32197
rect 13139 32373 13197 32385
rect 13139 32197 13151 32373
rect 13185 32197 13197 32373
rect 13139 32185 13197 32197
rect 13397 32373 13455 32385
rect 13397 32197 13409 32373
rect 13443 32197 13455 32373
rect 13397 32185 13455 32197
rect 25613 32297 25671 32309
rect 25613 32121 25625 32297
rect 25659 32121 25671 32297
rect 25613 32109 25671 32121
rect 25871 32297 25929 32309
rect 25871 32121 25883 32297
rect 25917 32121 25929 32297
rect 25871 32109 25929 32121
rect 26129 32297 26187 32309
rect 26129 32121 26141 32297
rect 26175 32121 26187 32297
rect 26129 32109 26187 32121
rect 7498 31172 7556 31184
rect 7498 30996 7510 31172
rect 7544 30996 7556 31172
rect 7498 30984 7556 30996
rect 7756 31172 7814 31184
rect 7756 30996 7768 31172
rect 7802 30996 7814 31172
rect 7756 30984 7814 30996
rect 8014 31172 8072 31184
rect 8014 30996 8026 31172
rect 8060 30996 8072 31172
rect 8014 30984 8072 30996
rect 8272 31172 8330 31184
rect 8272 30996 8284 31172
rect 8318 30996 8330 31172
rect 8272 30984 8330 30996
rect 8530 31172 8588 31184
rect 8530 30996 8542 31172
rect 8576 30996 8588 31172
rect 8530 30984 8588 30996
rect 8788 31172 8846 31184
rect 8788 30996 8800 31172
rect 8834 30996 8846 31172
rect 8788 30984 8846 30996
rect 9046 31172 9104 31184
rect 9046 30996 9058 31172
rect 9092 30996 9104 31172
rect 9046 30984 9104 30996
rect 9304 31172 9362 31184
rect 9304 30996 9316 31172
rect 9350 30996 9362 31172
rect 9304 30984 9362 30996
rect 9562 31172 9620 31184
rect 9562 30996 9574 31172
rect 9608 30996 9620 31172
rect 9562 30984 9620 30996
rect 9820 31172 9878 31184
rect 9820 30996 9832 31172
rect 9866 30996 9878 31172
rect 9820 30984 9878 30996
rect 10078 31172 10136 31184
rect 10078 30996 10090 31172
rect 10124 30996 10136 31172
rect 10078 30984 10136 30996
rect 10336 31172 10394 31184
rect 10336 30996 10348 31172
rect 10382 30996 10394 31172
rect 10336 30984 10394 30996
rect 10594 31172 10652 31184
rect 10594 30996 10606 31172
rect 10640 30996 10652 31172
rect 10594 30984 10652 30996
rect 12881 30913 12939 30925
rect 12881 30737 12893 30913
rect 12927 30737 12939 30913
rect 12881 30725 12939 30737
rect 13139 30913 13197 30925
rect 13139 30737 13151 30913
rect 13185 30737 13197 30913
rect 13139 30725 13197 30737
rect 13397 30913 13455 30925
rect 13397 30737 13409 30913
rect 13443 30737 13455 30913
rect 13397 30725 13455 30737
rect 12634 29465 12686 29477
rect 12634 29431 12642 29465
rect 12676 29431 12686 29465
rect 12634 29397 12686 29431
rect 12634 29363 12642 29397
rect 12676 29363 12686 29397
rect 12634 29277 12686 29363
rect 12716 29465 12770 29477
rect 12716 29431 12726 29465
rect 12760 29431 12770 29465
rect 12716 29397 12770 29431
rect 12716 29363 12726 29397
rect 12760 29363 12770 29397
rect 12716 29329 12770 29363
rect 12716 29295 12726 29329
rect 12760 29295 12770 29329
rect 12716 29277 12770 29295
rect 12800 29465 12854 29477
rect 12800 29431 12810 29465
rect 12844 29431 12854 29465
rect 12800 29397 12854 29431
rect 12800 29363 12810 29397
rect 12844 29363 12854 29397
rect 12800 29277 12854 29363
rect 12884 29465 12938 29477
rect 12884 29431 12894 29465
rect 12928 29431 12938 29465
rect 12884 29397 12938 29431
rect 12884 29363 12894 29397
rect 12928 29363 12938 29397
rect 12884 29329 12938 29363
rect 12884 29295 12894 29329
rect 12928 29295 12938 29329
rect 12884 29277 12938 29295
rect 12968 29465 13022 29477
rect 12968 29431 12978 29465
rect 13012 29431 13022 29465
rect 12968 29397 13022 29431
rect 12968 29363 12978 29397
rect 13012 29363 13022 29397
rect 12968 29277 13022 29363
rect 13052 29465 13106 29477
rect 13052 29431 13062 29465
rect 13096 29431 13106 29465
rect 13052 29397 13106 29431
rect 13052 29363 13062 29397
rect 13096 29363 13106 29397
rect 13052 29329 13106 29363
rect 13052 29295 13062 29329
rect 13096 29295 13106 29329
rect 13052 29277 13106 29295
rect 13136 29465 13190 29477
rect 13136 29431 13146 29465
rect 13180 29431 13190 29465
rect 13136 29397 13190 29431
rect 13136 29363 13146 29397
rect 13180 29363 13190 29397
rect 13136 29277 13190 29363
rect 13220 29465 13274 29477
rect 13220 29431 13230 29465
rect 13264 29431 13274 29465
rect 13220 29397 13274 29431
rect 13220 29363 13230 29397
rect 13264 29363 13274 29397
rect 13220 29329 13274 29363
rect 13220 29295 13230 29329
rect 13264 29295 13274 29329
rect 13220 29277 13274 29295
rect 13304 29465 13356 29477
rect 13304 29431 13314 29465
rect 13348 29431 13356 29465
rect 13304 29397 13356 29431
rect 13304 29363 13314 29397
rect 13348 29363 13356 29397
rect 13304 29277 13356 29363
rect 20230 31096 20288 31108
rect 20230 30920 20242 31096
rect 20276 30920 20288 31096
rect 20230 30908 20288 30920
rect 20488 31096 20546 31108
rect 20488 30920 20500 31096
rect 20534 30920 20546 31096
rect 20488 30908 20546 30920
rect 20746 31096 20804 31108
rect 20746 30920 20758 31096
rect 20792 30920 20804 31096
rect 20746 30908 20804 30920
rect 21004 31096 21062 31108
rect 21004 30920 21016 31096
rect 21050 30920 21062 31096
rect 21004 30908 21062 30920
rect 21262 31096 21320 31108
rect 21262 30920 21274 31096
rect 21308 30920 21320 31096
rect 21262 30908 21320 30920
rect 21520 31096 21578 31108
rect 21520 30920 21532 31096
rect 21566 30920 21578 31096
rect 21520 30908 21578 30920
rect 21778 31096 21836 31108
rect 21778 30920 21790 31096
rect 21824 30920 21836 31096
rect 21778 30908 21836 30920
rect 22036 31096 22094 31108
rect 22036 30920 22048 31096
rect 22082 30920 22094 31096
rect 22036 30908 22094 30920
rect 22294 31096 22352 31108
rect 22294 30920 22306 31096
rect 22340 30920 22352 31096
rect 22294 30908 22352 30920
rect 22552 31096 22610 31108
rect 22552 30920 22564 31096
rect 22598 30920 22610 31096
rect 22552 30908 22610 30920
rect 22810 31096 22868 31108
rect 22810 30920 22822 31096
rect 22856 30920 22868 31096
rect 22810 30908 22868 30920
rect 23068 31096 23126 31108
rect 23068 30920 23080 31096
rect 23114 30920 23126 31096
rect 23068 30908 23126 30920
rect 23326 31096 23384 31108
rect 23326 30920 23338 31096
rect 23372 30920 23384 31096
rect 23326 30908 23384 30920
rect 25613 30837 25671 30849
rect 25613 30661 25625 30837
rect 25659 30661 25671 30837
rect 25613 30649 25671 30661
rect 25871 30837 25929 30849
rect 25871 30661 25883 30837
rect 25917 30661 25929 30837
rect 25871 30649 25929 30661
rect 26129 30837 26187 30849
rect 26129 30661 26141 30837
rect 26175 30661 26187 30837
rect 26129 30649 26187 30661
rect 25366 29389 25418 29401
rect 25366 29355 25374 29389
rect 25408 29355 25418 29389
rect 25366 29321 25418 29355
rect 25366 29287 25374 29321
rect 25408 29287 25418 29321
rect 25366 29201 25418 29287
rect 25448 29389 25502 29401
rect 25448 29355 25458 29389
rect 25492 29355 25502 29389
rect 25448 29321 25502 29355
rect 25448 29287 25458 29321
rect 25492 29287 25502 29321
rect 25448 29253 25502 29287
rect 25448 29219 25458 29253
rect 25492 29219 25502 29253
rect 25448 29201 25502 29219
rect 25532 29389 25586 29401
rect 25532 29355 25542 29389
rect 25576 29355 25586 29389
rect 25532 29321 25586 29355
rect 25532 29287 25542 29321
rect 25576 29287 25586 29321
rect 25532 29201 25586 29287
rect 25616 29389 25670 29401
rect 25616 29355 25626 29389
rect 25660 29355 25670 29389
rect 25616 29321 25670 29355
rect 25616 29287 25626 29321
rect 25660 29287 25670 29321
rect 25616 29253 25670 29287
rect 25616 29219 25626 29253
rect 25660 29219 25670 29253
rect 25616 29201 25670 29219
rect 25700 29389 25754 29401
rect 25700 29355 25710 29389
rect 25744 29355 25754 29389
rect 25700 29321 25754 29355
rect 25700 29287 25710 29321
rect 25744 29287 25754 29321
rect 25700 29201 25754 29287
rect 25784 29389 25838 29401
rect 25784 29355 25794 29389
rect 25828 29355 25838 29389
rect 25784 29321 25838 29355
rect 25784 29287 25794 29321
rect 25828 29287 25838 29321
rect 25784 29253 25838 29287
rect 25784 29219 25794 29253
rect 25828 29219 25838 29253
rect 25784 29201 25838 29219
rect 25868 29389 25922 29401
rect 25868 29355 25878 29389
rect 25912 29355 25922 29389
rect 25868 29321 25922 29355
rect 25868 29287 25878 29321
rect 25912 29287 25922 29321
rect 25868 29201 25922 29287
rect 25952 29389 26006 29401
rect 25952 29355 25962 29389
rect 25996 29355 26006 29389
rect 25952 29321 26006 29355
rect 25952 29287 25962 29321
rect 25996 29287 26006 29321
rect 25952 29253 26006 29287
rect 25952 29219 25962 29253
rect 25996 29219 26006 29253
rect 25952 29201 26006 29219
rect 26036 29389 26088 29401
rect 26036 29355 26046 29389
rect 26080 29355 26088 29389
rect 26036 29321 26088 29355
rect 26036 29287 26046 29321
rect 26080 29287 26088 29321
rect 26036 29201 26088 29287
rect 13001 25669 13059 25681
rect 13001 25493 13013 25669
rect 13047 25493 13059 25669
rect 13001 25481 13059 25493
rect 13259 25669 13317 25681
rect 13259 25493 13271 25669
rect 13305 25493 13317 25669
rect 13259 25481 13317 25493
rect 13517 25669 13575 25681
rect 13517 25493 13529 25669
rect 13563 25493 13575 25669
rect 13517 25481 13575 25493
rect 25709 25539 25767 25551
rect 25709 25363 25721 25539
rect 25755 25363 25767 25539
rect 25709 25351 25767 25363
rect 25967 25539 26025 25551
rect 25967 25363 25979 25539
rect 26013 25363 26025 25539
rect 25967 25351 26025 25363
rect 26225 25539 26283 25551
rect 26225 25363 26237 25539
rect 26271 25363 26283 25539
rect 26225 25351 26283 25363
rect 7618 24468 7676 24480
rect 7618 24292 7630 24468
rect 7664 24292 7676 24468
rect 7618 24280 7676 24292
rect 7876 24468 7934 24480
rect 7876 24292 7888 24468
rect 7922 24292 7934 24468
rect 7876 24280 7934 24292
rect 8134 24468 8192 24480
rect 8134 24292 8146 24468
rect 8180 24292 8192 24468
rect 8134 24280 8192 24292
rect 8392 24468 8450 24480
rect 8392 24292 8404 24468
rect 8438 24292 8450 24468
rect 8392 24280 8450 24292
rect 8650 24468 8708 24480
rect 8650 24292 8662 24468
rect 8696 24292 8708 24468
rect 8650 24280 8708 24292
rect 8908 24468 8966 24480
rect 8908 24292 8920 24468
rect 8954 24292 8966 24468
rect 8908 24280 8966 24292
rect 9166 24468 9224 24480
rect 9166 24292 9178 24468
rect 9212 24292 9224 24468
rect 9166 24280 9224 24292
rect 9424 24468 9482 24480
rect 9424 24292 9436 24468
rect 9470 24292 9482 24468
rect 9424 24280 9482 24292
rect 9682 24468 9740 24480
rect 9682 24292 9694 24468
rect 9728 24292 9740 24468
rect 9682 24280 9740 24292
rect 9940 24468 9998 24480
rect 9940 24292 9952 24468
rect 9986 24292 9998 24468
rect 9940 24280 9998 24292
rect 10198 24468 10256 24480
rect 10198 24292 10210 24468
rect 10244 24292 10256 24468
rect 10198 24280 10256 24292
rect 10456 24468 10514 24480
rect 10456 24292 10468 24468
rect 10502 24292 10514 24468
rect 10456 24280 10514 24292
rect 10714 24468 10772 24480
rect 10714 24292 10726 24468
rect 10760 24292 10772 24468
rect 10714 24280 10772 24292
rect 13001 24209 13059 24221
rect 13001 24033 13013 24209
rect 13047 24033 13059 24209
rect 13001 24021 13059 24033
rect 13259 24209 13317 24221
rect 13259 24033 13271 24209
rect 13305 24033 13317 24209
rect 13259 24021 13317 24033
rect 13517 24209 13575 24221
rect 13517 24033 13529 24209
rect 13563 24033 13575 24209
rect 13517 24021 13575 24033
rect 12754 22761 12806 22773
rect 12754 22727 12762 22761
rect 12796 22727 12806 22761
rect 12754 22693 12806 22727
rect 12754 22659 12762 22693
rect 12796 22659 12806 22693
rect 12754 22573 12806 22659
rect 12836 22761 12890 22773
rect 12836 22727 12846 22761
rect 12880 22727 12890 22761
rect 12836 22693 12890 22727
rect 12836 22659 12846 22693
rect 12880 22659 12890 22693
rect 12836 22625 12890 22659
rect 12836 22591 12846 22625
rect 12880 22591 12890 22625
rect 12836 22573 12890 22591
rect 12920 22761 12974 22773
rect 12920 22727 12930 22761
rect 12964 22727 12974 22761
rect 12920 22693 12974 22727
rect 12920 22659 12930 22693
rect 12964 22659 12974 22693
rect 12920 22573 12974 22659
rect 13004 22761 13058 22773
rect 13004 22727 13014 22761
rect 13048 22727 13058 22761
rect 13004 22693 13058 22727
rect 13004 22659 13014 22693
rect 13048 22659 13058 22693
rect 13004 22625 13058 22659
rect 13004 22591 13014 22625
rect 13048 22591 13058 22625
rect 13004 22573 13058 22591
rect 13088 22761 13142 22773
rect 13088 22727 13098 22761
rect 13132 22727 13142 22761
rect 13088 22693 13142 22727
rect 13088 22659 13098 22693
rect 13132 22659 13142 22693
rect 13088 22573 13142 22659
rect 13172 22761 13226 22773
rect 13172 22727 13182 22761
rect 13216 22727 13226 22761
rect 13172 22693 13226 22727
rect 13172 22659 13182 22693
rect 13216 22659 13226 22693
rect 13172 22625 13226 22659
rect 13172 22591 13182 22625
rect 13216 22591 13226 22625
rect 13172 22573 13226 22591
rect 13256 22761 13310 22773
rect 13256 22727 13266 22761
rect 13300 22727 13310 22761
rect 13256 22693 13310 22727
rect 13256 22659 13266 22693
rect 13300 22659 13310 22693
rect 13256 22573 13310 22659
rect 13340 22761 13394 22773
rect 13340 22727 13350 22761
rect 13384 22727 13394 22761
rect 13340 22693 13394 22727
rect 13340 22659 13350 22693
rect 13384 22659 13394 22693
rect 13340 22625 13394 22659
rect 13340 22591 13350 22625
rect 13384 22591 13394 22625
rect 13340 22573 13394 22591
rect 13424 22761 13476 22773
rect 13424 22727 13434 22761
rect 13468 22727 13476 22761
rect 13424 22693 13476 22727
rect 13424 22659 13434 22693
rect 13468 22659 13476 22693
rect 13424 22573 13476 22659
rect 20326 24338 20384 24350
rect 20326 24162 20338 24338
rect 20372 24162 20384 24338
rect 20326 24150 20384 24162
rect 20584 24338 20642 24350
rect 20584 24162 20596 24338
rect 20630 24162 20642 24338
rect 20584 24150 20642 24162
rect 20842 24338 20900 24350
rect 20842 24162 20854 24338
rect 20888 24162 20900 24338
rect 20842 24150 20900 24162
rect 21100 24338 21158 24350
rect 21100 24162 21112 24338
rect 21146 24162 21158 24338
rect 21100 24150 21158 24162
rect 21358 24338 21416 24350
rect 21358 24162 21370 24338
rect 21404 24162 21416 24338
rect 21358 24150 21416 24162
rect 21616 24338 21674 24350
rect 21616 24162 21628 24338
rect 21662 24162 21674 24338
rect 21616 24150 21674 24162
rect 21874 24338 21932 24350
rect 21874 24162 21886 24338
rect 21920 24162 21932 24338
rect 21874 24150 21932 24162
rect 22132 24338 22190 24350
rect 22132 24162 22144 24338
rect 22178 24162 22190 24338
rect 22132 24150 22190 24162
rect 22390 24338 22448 24350
rect 22390 24162 22402 24338
rect 22436 24162 22448 24338
rect 22390 24150 22448 24162
rect 22648 24338 22706 24350
rect 22648 24162 22660 24338
rect 22694 24162 22706 24338
rect 22648 24150 22706 24162
rect 22906 24338 22964 24350
rect 22906 24162 22918 24338
rect 22952 24162 22964 24338
rect 22906 24150 22964 24162
rect 23164 24338 23222 24350
rect 23164 24162 23176 24338
rect 23210 24162 23222 24338
rect 23164 24150 23222 24162
rect 23422 24338 23480 24350
rect 23422 24162 23434 24338
rect 23468 24162 23480 24338
rect 23422 24150 23480 24162
rect 25709 24079 25767 24091
rect 25709 23903 25721 24079
rect 25755 23903 25767 24079
rect 25709 23891 25767 23903
rect 25967 24079 26025 24091
rect 25967 23903 25979 24079
rect 26013 23903 26025 24079
rect 25967 23891 26025 23903
rect 26225 24079 26283 24091
rect 26225 23903 26237 24079
rect 26271 23903 26283 24079
rect 26225 23891 26283 23903
rect 25462 22631 25514 22643
rect 25462 22597 25470 22631
rect 25504 22597 25514 22631
rect 25462 22563 25514 22597
rect 25462 22529 25470 22563
rect 25504 22529 25514 22563
rect 25462 22443 25514 22529
rect 25544 22631 25598 22643
rect 25544 22597 25554 22631
rect 25588 22597 25598 22631
rect 25544 22563 25598 22597
rect 25544 22529 25554 22563
rect 25588 22529 25598 22563
rect 25544 22495 25598 22529
rect 25544 22461 25554 22495
rect 25588 22461 25598 22495
rect 25544 22443 25598 22461
rect 25628 22631 25682 22643
rect 25628 22597 25638 22631
rect 25672 22597 25682 22631
rect 25628 22563 25682 22597
rect 25628 22529 25638 22563
rect 25672 22529 25682 22563
rect 25628 22443 25682 22529
rect 25712 22631 25766 22643
rect 25712 22597 25722 22631
rect 25756 22597 25766 22631
rect 25712 22563 25766 22597
rect 25712 22529 25722 22563
rect 25756 22529 25766 22563
rect 25712 22495 25766 22529
rect 25712 22461 25722 22495
rect 25756 22461 25766 22495
rect 25712 22443 25766 22461
rect 25796 22631 25850 22643
rect 25796 22597 25806 22631
rect 25840 22597 25850 22631
rect 25796 22563 25850 22597
rect 25796 22529 25806 22563
rect 25840 22529 25850 22563
rect 25796 22443 25850 22529
rect 25880 22631 25934 22643
rect 25880 22597 25890 22631
rect 25924 22597 25934 22631
rect 25880 22563 25934 22597
rect 25880 22529 25890 22563
rect 25924 22529 25934 22563
rect 25880 22495 25934 22529
rect 25880 22461 25890 22495
rect 25924 22461 25934 22495
rect 25880 22443 25934 22461
rect 25964 22631 26018 22643
rect 25964 22597 25974 22631
rect 26008 22597 26018 22631
rect 25964 22563 26018 22597
rect 25964 22529 25974 22563
rect 26008 22529 26018 22563
rect 25964 22443 26018 22529
rect 26048 22631 26102 22643
rect 26048 22597 26058 22631
rect 26092 22597 26102 22631
rect 26048 22563 26102 22597
rect 26048 22529 26058 22563
rect 26092 22529 26102 22563
rect 26048 22495 26102 22529
rect 26048 22461 26058 22495
rect 26092 22461 26102 22495
rect 26048 22443 26102 22461
rect 26132 22631 26184 22643
rect 26132 22597 26142 22631
rect 26176 22597 26184 22631
rect 26132 22563 26184 22597
rect 26132 22529 26142 22563
rect 26176 22529 26184 22563
rect 26132 22443 26184 22529
rect 12877 18623 12935 18635
rect 12877 18447 12889 18623
rect 12923 18447 12935 18623
rect 12877 18435 12935 18447
rect 13135 18623 13193 18635
rect 13135 18447 13147 18623
rect 13181 18447 13193 18623
rect 13135 18435 13193 18447
rect 13393 18623 13451 18635
rect 13393 18447 13405 18623
rect 13439 18447 13451 18623
rect 13393 18435 13451 18447
rect 26059 18493 26117 18505
rect 26059 18317 26071 18493
rect 26105 18317 26117 18493
rect 26059 18305 26117 18317
rect 26317 18493 26375 18505
rect 26317 18317 26329 18493
rect 26363 18317 26375 18493
rect 26317 18305 26375 18317
rect 26575 18493 26633 18505
rect 26575 18317 26587 18493
rect 26621 18317 26633 18493
rect 26575 18305 26633 18317
rect 7494 17422 7552 17434
rect 7494 17246 7506 17422
rect 7540 17246 7552 17422
rect 7494 17234 7552 17246
rect 7752 17422 7810 17434
rect 7752 17246 7764 17422
rect 7798 17246 7810 17422
rect 7752 17234 7810 17246
rect 8010 17422 8068 17434
rect 8010 17246 8022 17422
rect 8056 17246 8068 17422
rect 8010 17234 8068 17246
rect 8268 17422 8326 17434
rect 8268 17246 8280 17422
rect 8314 17246 8326 17422
rect 8268 17234 8326 17246
rect 8526 17422 8584 17434
rect 8526 17246 8538 17422
rect 8572 17246 8584 17422
rect 8526 17234 8584 17246
rect 8784 17422 8842 17434
rect 8784 17246 8796 17422
rect 8830 17246 8842 17422
rect 8784 17234 8842 17246
rect 9042 17422 9100 17434
rect 9042 17246 9054 17422
rect 9088 17246 9100 17422
rect 9042 17234 9100 17246
rect 9300 17422 9358 17434
rect 9300 17246 9312 17422
rect 9346 17246 9358 17422
rect 9300 17234 9358 17246
rect 9558 17422 9616 17434
rect 9558 17246 9570 17422
rect 9604 17246 9616 17422
rect 9558 17234 9616 17246
rect 9816 17422 9874 17434
rect 9816 17246 9828 17422
rect 9862 17246 9874 17422
rect 9816 17234 9874 17246
rect 10074 17422 10132 17434
rect 10074 17246 10086 17422
rect 10120 17246 10132 17422
rect 10074 17234 10132 17246
rect 10332 17422 10390 17434
rect 10332 17246 10344 17422
rect 10378 17246 10390 17422
rect 10332 17234 10390 17246
rect 10590 17422 10648 17434
rect 10590 17246 10602 17422
rect 10636 17246 10648 17422
rect 10590 17234 10648 17246
rect 12877 17163 12935 17175
rect 12877 16987 12889 17163
rect 12923 16987 12935 17163
rect 12877 16975 12935 16987
rect 13135 17163 13193 17175
rect 13135 16987 13147 17163
rect 13181 16987 13193 17163
rect 13135 16975 13193 16987
rect 13393 17163 13451 17175
rect 13393 16987 13405 17163
rect 13439 16987 13451 17163
rect 13393 16975 13451 16987
rect 12630 15715 12682 15727
rect 12630 15681 12638 15715
rect 12672 15681 12682 15715
rect 12630 15647 12682 15681
rect 12630 15613 12638 15647
rect 12672 15613 12682 15647
rect 12630 15527 12682 15613
rect 12712 15715 12766 15727
rect 12712 15681 12722 15715
rect 12756 15681 12766 15715
rect 12712 15647 12766 15681
rect 12712 15613 12722 15647
rect 12756 15613 12766 15647
rect 12712 15579 12766 15613
rect 12712 15545 12722 15579
rect 12756 15545 12766 15579
rect 12712 15527 12766 15545
rect 12796 15715 12850 15727
rect 12796 15681 12806 15715
rect 12840 15681 12850 15715
rect 12796 15647 12850 15681
rect 12796 15613 12806 15647
rect 12840 15613 12850 15647
rect 12796 15527 12850 15613
rect 12880 15715 12934 15727
rect 12880 15681 12890 15715
rect 12924 15681 12934 15715
rect 12880 15647 12934 15681
rect 12880 15613 12890 15647
rect 12924 15613 12934 15647
rect 12880 15579 12934 15613
rect 12880 15545 12890 15579
rect 12924 15545 12934 15579
rect 12880 15527 12934 15545
rect 12964 15715 13018 15727
rect 12964 15681 12974 15715
rect 13008 15681 13018 15715
rect 12964 15647 13018 15681
rect 12964 15613 12974 15647
rect 13008 15613 13018 15647
rect 12964 15527 13018 15613
rect 13048 15715 13102 15727
rect 13048 15681 13058 15715
rect 13092 15681 13102 15715
rect 13048 15647 13102 15681
rect 13048 15613 13058 15647
rect 13092 15613 13102 15647
rect 13048 15579 13102 15613
rect 13048 15545 13058 15579
rect 13092 15545 13102 15579
rect 13048 15527 13102 15545
rect 13132 15715 13186 15727
rect 13132 15681 13142 15715
rect 13176 15681 13186 15715
rect 13132 15647 13186 15681
rect 13132 15613 13142 15647
rect 13176 15613 13186 15647
rect 13132 15527 13186 15613
rect 13216 15715 13270 15727
rect 13216 15681 13226 15715
rect 13260 15681 13270 15715
rect 13216 15647 13270 15681
rect 13216 15613 13226 15647
rect 13260 15613 13270 15647
rect 13216 15579 13270 15613
rect 13216 15545 13226 15579
rect 13260 15545 13270 15579
rect 13216 15527 13270 15545
rect 13300 15715 13352 15727
rect 13300 15681 13310 15715
rect 13344 15681 13352 15715
rect 13300 15647 13352 15681
rect 13300 15613 13310 15647
rect 13344 15613 13352 15647
rect 13300 15527 13352 15613
rect 20676 17292 20734 17304
rect 20676 17116 20688 17292
rect 20722 17116 20734 17292
rect 20676 17104 20734 17116
rect 20934 17292 20992 17304
rect 20934 17116 20946 17292
rect 20980 17116 20992 17292
rect 20934 17104 20992 17116
rect 21192 17292 21250 17304
rect 21192 17116 21204 17292
rect 21238 17116 21250 17292
rect 21192 17104 21250 17116
rect 21450 17292 21508 17304
rect 21450 17116 21462 17292
rect 21496 17116 21508 17292
rect 21450 17104 21508 17116
rect 21708 17292 21766 17304
rect 21708 17116 21720 17292
rect 21754 17116 21766 17292
rect 21708 17104 21766 17116
rect 21966 17292 22024 17304
rect 21966 17116 21978 17292
rect 22012 17116 22024 17292
rect 21966 17104 22024 17116
rect 22224 17292 22282 17304
rect 22224 17116 22236 17292
rect 22270 17116 22282 17292
rect 22224 17104 22282 17116
rect 22482 17292 22540 17304
rect 22482 17116 22494 17292
rect 22528 17116 22540 17292
rect 22482 17104 22540 17116
rect 22740 17292 22798 17304
rect 22740 17116 22752 17292
rect 22786 17116 22798 17292
rect 22740 17104 22798 17116
rect 22998 17292 23056 17304
rect 22998 17116 23010 17292
rect 23044 17116 23056 17292
rect 22998 17104 23056 17116
rect 23256 17292 23314 17304
rect 23256 17116 23268 17292
rect 23302 17116 23314 17292
rect 23256 17104 23314 17116
rect 23514 17292 23572 17304
rect 23514 17116 23526 17292
rect 23560 17116 23572 17292
rect 23514 17104 23572 17116
rect 23772 17292 23830 17304
rect 23772 17116 23784 17292
rect 23818 17116 23830 17292
rect 23772 17104 23830 17116
rect 26059 17033 26117 17045
rect 26059 16857 26071 17033
rect 26105 16857 26117 17033
rect 26059 16845 26117 16857
rect 26317 17033 26375 17045
rect 26317 16857 26329 17033
rect 26363 16857 26375 17033
rect 26317 16845 26375 16857
rect 26575 17033 26633 17045
rect 26575 16857 26587 17033
rect 26621 16857 26633 17033
rect 26575 16845 26633 16857
rect 25812 15585 25864 15597
rect 25812 15551 25820 15585
rect 25854 15551 25864 15585
rect 25812 15517 25864 15551
rect 25812 15483 25820 15517
rect 25854 15483 25864 15517
rect 25812 15397 25864 15483
rect 25894 15585 25948 15597
rect 25894 15551 25904 15585
rect 25938 15551 25948 15585
rect 25894 15517 25948 15551
rect 25894 15483 25904 15517
rect 25938 15483 25948 15517
rect 25894 15449 25948 15483
rect 25894 15415 25904 15449
rect 25938 15415 25948 15449
rect 25894 15397 25948 15415
rect 25978 15585 26032 15597
rect 25978 15551 25988 15585
rect 26022 15551 26032 15585
rect 25978 15517 26032 15551
rect 25978 15483 25988 15517
rect 26022 15483 26032 15517
rect 25978 15397 26032 15483
rect 26062 15585 26116 15597
rect 26062 15551 26072 15585
rect 26106 15551 26116 15585
rect 26062 15517 26116 15551
rect 26062 15483 26072 15517
rect 26106 15483 26116 15517
rect 26062 15449 26116 15483
rect 26062 15415 26072 15449
rect 26106 15415 26116 15449
rect 26062 15397 26116 15415
rect 26146 15585 26200 15597
rect 26146 15551 26156 15585
rect 26190 15551 26200 15585
rect 26146 15517 26200 15551
rect 26146 15483 26156 15517
rect 26190 15483 26200 15517
rect 26146 15397 26200 15483
rect 26230 15585 26284 15597
rect 26230 15551 26240 15585
rect 26274 15551 26284 15585
rect 26230 15517 26284 15551
rect 26230 15483 26240 15517
rect 26274 15483 26284 15517
rect 26230 15449 26284 15483
rect 26230 15415 26240 15449
rect 26274 15415 26284 15449
rect 26230 15397 26284 15415
rect 26314 15585 26368 15597
rect 26314 15551 26324 15585
rect 26358 15551 26368 15585
rect 26314 15517 26368 15551
rect 26314 15483 26324 15517
rect 26358 15483 26368 15517
rect 26314 15397 26368 15483
rect 26398 15585 26452 15597
rect 26398 15551 26408 15585
rect 26442 15551 26452 15585
rect 26398 15517 26452 15551
rect 26398 15483 26408 15517
rect 26442 15483 26452 15517
rect 26398 15449 26452 15483
rect 26398 15415 26408 15449
rect 26442 15415 26452 15449
rect 26398 15397 26452 15415
rect 26482 15585 26534 15597
rect 26482 15551 26492 15585
rect 26526 15551 26534 15585
rect 26482 15517 26534 15551
rect 26482 15483 26492 15517
rect 26526 15483 26534 15517
rect 26482 15397 26534 15483
<< ndiffc >>
rect 7490 36495 7524 36671
rect 7748 36495 7782 36671
rect 8006 36495 8040 36671
rect 8264 36495 8298 36671
rect 8522 36495 8556 36671
rect 8780 36495 8814 36671
rect 9038 36495 9072 36671
rect 9296 36495 9330 36671
rect 9554 36495 9588 36671
rect 9812 36495 9846 36671
rect 10070 36495 10104 36671
rect 10328 36495 10362 36671
rect 10586 36495 10620 36671
rect 7490 36175 7524 36235
rect 7748 36175 7782 36235
rect 8006 36175 8040 36235
rect 8264 36175 8298 36235
rect 8522 36175 8556 36235
rect 8780 36175 8814 36235
rect 9038 36175 9072 36235
rect 9296 36175 9330 36235
rect 9554 36175 9588 36235
rect 9812 36175 9846 36235
rect 10070 36175 10104 36235
rect 10328 36175 10362 36235
rect 10586 36175 10620 36235
rect 12873 37627 12907 37803
rect 13131 37627 13165 37803
rect 13389 37627 13423 37803
rect 12873 36167 12907 36343
rect 13131 36167 13165 36343
rect 13389 36167 13423 36343
rect 20278 36613 20312 36789
rect 20536 36613 20570 36789
rect 20794 36613 20828 36789
rect 21052 36613 21086 36789
rect 21310 36613 21344 36789
rect 21568 36613 21602 36789
rect 21826 36613 21860 36789
rect 22084 36613 22118 36789
rect 22342 36613 22376 36789
rect 22600 36613 22634 36789
rect 22858 36613 22892 36789
rect 23116 36613 23150 36789
rect 23374 36613 23408 36789
rect 20278 36293 20312 36353
rect 20536 36293 20570 36353
rect 20794 36293 20828 36353
rect 21052 36293 21086 36353
rect 21310 36293 21344 36353
rect 21568 36293 21602 36353
rect 21826 36293 21860 36353
rect 22084 36293 22118 36353
rect 22342 36293 22376 36353
rect 22600 36293 22634 36353
rect 22858 36293 22892 36353
rect 23116 36293 23150 36353
rect 23374 36293 23408 36353
rect 12622 34965 12656 34999
rect 12706 35033 12740 35067
rect 12706 34965 12740 34999
rect 12790 34965 12824 34999
rect 12874 35033 12908 35067
rect 12874 34965 12908 34999
rect 12958 34965 12992 34999
rect 13042 35033 13076 35067
rect 13042 34965 13076 34999
rect 13126 34965 13160 34999
rect 13210 35033 13244 35067
rect 13210 34965 13244 34999
rect 13294 34965 13328 34999
rect 25661 37745 25695 37921
rect 25919 37745 25953 37921
rect 26177 37745 26211 37921
rect 25661 36285 25695 36461
rect 25919 36285 25953 36461
rect 26177 36285 26211 36461
rect 25410 35083 25444 35117
rect 25494 35151 25528 35185
rect 25494 35083 25528 35117
rect 25578 35083 25612 35117
rect 25662 35151 25696 35185
rect 25662 35083 25696 35117
rect 25746 35083 25780 35117
rect 25830 35151 25864 35185
rect 25830 35083 25864 35117
rect 25914 35083 25948 35117
rect 25998 35151 26032 35185
rect 25998 35083 26032 35117
rect 26082 35083 26116 35117
rect 7510 30569 7544 30745
rect 7768 30569 7802 30745
rect 8026 30569 8060 30745
rect 8284 30569 8318 30745
rect 8542 30569 8576 30745
rect 8800 30569 8834 30745
rect 9058 30569 9092 30745
rect 9316 30569 9350 30745
rect 9574 30569 9608 30745
rect 9832 30569 9866 30745
rect 10090 30569 10124 30745
rect 10348 30569 10382 30745
rect 10606 30569 10640 30745
rect 7510 30249 7544 30309
rect 7768 30249 7802 30309
rect 8026 30249 8060 30309
rect 8284 30249 8318 30309
rect 8542 30249 8576 30309
rect 8800 30249 8834 30309
rect 9058 30249 9092 30309
rect 9316 30249 9350 30309
rect 9574 30249 9608 30309
rect 9832 30249 9866 30309
rect 10090 30249 10124 30309
rect 10348 30249 10382 30309
rect 10606 30249 10640 30309
rect 12893 31701 12927 31877
rect 13151 31701 13185 31877
rect 13409 31701 13443 31877
rect 12893 30241 12927 30417
rect 13151 30241 13185 30417
rect 13409 30241 13443 30417
rect 20242 30493 20276 30669
rect 20500 30493 20534 30669
rect 20758 30493 20792 30669
rect 21016 30493 21050 30669
rect 21274 30493 21308 30669
rect 21532 30493 21566 30669
rect 21790 30493 21824 30669
rect 22048 30493 22082 30669
rect 22306 30493 22340 30669
rect 22564 30493 22598 30669
rect 22822 30493 22856 30669
rect 23080 30493 23114 30669
rect 23338 30493 23372 30669
rect 20242 30173 20276 30233
rect 20500 30173 20534 30233
rect 20758 30173 20792 30233
rect 21016 30173 21050 30233
rect 21274 30173 21308 30233
rect 21532 30173 21566 30233
rect 21790 30173 21824 30233
rect 22048 30173 22082 30233
rect 22306 30173 22340 30233
rect 22564 30173 22598 30233
rect 22822 30173 22856 30233
rect 23080 30173 23114 30233
rect 23338 30173 23372 30233
rect 12642 29039 12676 29073
rect 12726 29107 12760 29141
rect 12726 29039 12760 29073
rect 12810 29039 12844 29073
rect 12894 29107 12928 29141
rect 12894 29039 12928 29073
rect 12978 29039 13012 29073
rect 13062 29107 13096 29141
rect 13062 29039 13096 29073
rect 13146 29039 13180 29073
rect 13230 29107 13264 29141
rect 13230 29039 13264 29073
rect 13314 29039 13348 29073
rect 25625 31625 25659 31801
rect 25883 31625 25917 31801
rect 26141 31625 26175 31801
rect 25625 30165 25659 30341
rect 25883 30165 25917 30341
rect 26141 30165 26175 30341
rect 25374 28963 25408 28997
rect 25458 29031 25492 29065
rect 25458 28963 25492 28997
rect 25542 28963 25576 28997
rect 25626 29031 25660 29065
rect 25626 28963 25660 28997
rect 25710 28963 25744 28997
rect 25794 29031 25828 29065
rect 25794 28963 25828 28997
rect 25878 28963 25912 28997
rect 25962 29031 25996 29065
rect 25962 28963 25996 28997
rect 26046 28963 26080 28997
rect 7630 23865 7664 24041
rect 7888 23865 7922 24041
rect 8146 23865 8180 24041
rect 8404 23865 8438 24041
rect 8662 23865 8696 24041
rect 8920 23865 8954 24041
rect 9178 23865 9212 24041
rect 9436 23865 9470 24041
rect 9694 23865 9728 24041
rect 9952 23865 9986 24041
rect 10210 23865 10244 24041
rect 10468 23865 10502 24041
rect 10726 23865 10760 24041
rect 7630 23545 7664 23605
rect 7888 23545 7922 23605
rect 8146 23545 8180 23605
rect 8404 23545 8438 23605
rect 8662 23545 8696 23605
rect 8920 23545 8954 23605
rect 9178 23545 9212 23605
rect 9436 23545 9470 23605
rect 9694 23545 9728 23605
rect 9952 23545 9986 23605
rect 10210 23545 10244 23605
rect 10468 23545 10502 23605
rect 10726 23545 10760 23605
rect 13013 24997 13047 25173
rect 13271 24997 13305 25173
rect 13529 24997 13563 25173
rect 13013 23537 13047 23713
rect 13271 23537 13305 23713
rect 13529 23537 13563 23713
rect 20338 23735 20372 23911
rect 20596 23735 20630 23911
rect 20854 23735 20888 23911
rect 21112 23735 21146 23911
rect 21370 23735 21404 23911
rect 21628 23735 21662 23911
rect 21886 23735 21920 23911
rect 22144 23735 22178 23911
rect 22402 23735 22436 23911
rect 22660 23735 22694 23911
rect 22918 23735 22952 23911
rect 23176 23735 23210 23911
rect 23434 23735 23468 23911
rect 20338 23415 20372 23475
rect 20596 23415 20630 23475
rect 20854 23415 20888 23475
rect 21112 23415 21146 23475
rect 21370 23415 21404 23475
rect 21628 23415 21662 23475
rect 21886 23415 21920 23475
rect 22144 23415 22178 23475
rect 22402 23415 22436 23475
rect 22660 23415 22694 23475
rect 22918 23415 22952 23475
rect 23176 23415 23210 23475
rect 23434 23415 23468 23475
rect 12762 22335 12796 22369
rect 12846 22403 12880 22437
rect 12846 22335 12880 22369
rect 12930 22335 12964 22369
rect 13014 22403 13048 22437
rect 13014 22335 13048 22369
rect 13098 22335 13132 22369
rect 13182 22403 13216 22437
rect 13182 22335 13216 22369
rect 13266 22335 13300 22369
rect 13350 22403 13384 22437
rect 13350 22335 13384 22369
rect 13434 22335 13468 22369
rect 25721 24867 25755 25043
rect 25979 24867 26013 25043
rect 26237 24867 26271 25043
rect 25721 23407 25755 23583
rect 25979 23407 26013 23583
rect 26237 23407 26271 23583
rect 25470 22205 25504 22239
rect 25554 22273 25588 22307
rect 25554 22205 25588 22239
rect 25638 22205 25672 22239
rect 25722 22273 25756 22307
rect 25722 22205 25756 22239
rect 25806 22205 25840 22239
rect 25890 22273 25924 22307
rect 25890 22205 25924 22239
rect 25974 22205 26008 22239
rect 26058 22273 26092 22307
rect 26058 22205 26092 22239
rect 26142 22205 26176 22239
rect 7506 16819 7540 16995
rect 7764 16819 7798 16995
rect 8022 16819 8056 16995
rect 8280 16819 8314 16995
rect 8538 16819 8572 16995
rect 8796 16819 8830 16995
rect 9054 16819 9088 16995
rect 9312 16819 9346 16995
rect 9570 16819 9604 16995
rect 9828 16819 9862 16995
rect 10086 16819 10120 16995
rect 10344 16819 10378 16995
rect 10602 16819 10636 16995
rect 7506 16499 7540 16559
rect 7764 16499 7798 16559
rect 8022 16499 8056 16559
rect 8280 16499 8314 16559
rect 8538 16499 8572 16559
rect 8796 16499 8830 16559
rect 9054 16499 9088 16559
rect 9312 16499 9346 16559
rect 9570 16499 9604 16559
rect 9828 16499 9862 16559
rect 10086 16499 10120 16559
rect 10344 16499 10378 16559
rect 10602 16499 10636 16559
rect 12889 17951 12923 18127
rect 13147 17951 13181 18127
rect 13405 17951 13439 18127
rect 12889 16491 12923 16667
rect 13147 16491 13181 16667
rect 13405 16491 13439 16667
rect 20688 16689 20722 16865
rect 20946 16689 20980 16865
rect 21204 16689 21238 16865
rect 21462 16689 21496 16865
rect 21720 16689 21754 16865
rect 21978 16689 22012 16865
rect 22236 16689 22270 16865
rect 22494 16689 22528 16865
rect 22752 16689 22786 16865
rect 23010 16689 23044 16865
rect 23268 16689 23302 16865
rect 23526 16689 23560 16865
rect 23784 16689 23818 16865
rect 20688 16369 20722 16429
rect 20946 16369 20980 16429
rect 21204 16369 21238 16429
rect 21462 16369 21496 16429
rect 21720 16369 21754 16429
rect 21978 16369 22012 16429
rect 22236 16369 22270 16429
rect 22494 16369 22528 16429
rect 22752 16369 22786 16429
rect 23010 16369 23044 16429
rect 23268 16369 23302 16429
rect 23526 16369 23560 16429
rect 23784 16369 23818 16429
rect 12638 15289 12672 15323
rect 12722 15357 12756 15391
rect 12722 15289 12756 15323
rect 12806 15289 12840 15323
rect 12890 15357 12924 15391
rect 12890 15289 12924 15323
rect 12974 15289 13008 15323
rect 13058 15357 13092 15391
rect 13058 15289 13092 15323
rect 13142 15289 13176 15323
rect 13226 15357 13260 15391
rect 13226 15289 13260 15323
rect 13310 15289 13344 15323
rect 26071 17821 26105 17997
rect 26329 17821 26363 17997
rect 26587 17821 26621 17997
rect 26071 16361 26105 16537
rect 26329 16361 26363 16537
rect 26587 16361 26621 16537
rect 25820 15159 25854 15193
rect 25904 15227 25938 15261
rect 25904 15159 25938 15193
rect 25988 15159 26022 15193
rect 26072 15227 26106 15261
rect 26072 15159 26106 15193
rect 26156 15159 26190 15193
rect 26240 15227 26274 15261
rect 26240 15159 26274 15193
rect 26324 15159 26358 15193
rect 26408 15227 26442 15261
rect 26408 15159 26442 15193
rect 26492 15159 26526 15193
<< pdiffc >>
rect 12873 38123 12907 38299
rect 13131 38123 13165 38299
rect 13389 38123 13423 38299
rect 25661 38241 25695 38417
rect 25919 38241 25953 38417
rect 26177 38241 26211 38417
rect 7490 36922 7524 37098
rect 7748 36922 7782 37098
rect 8006 36922 8040 37098
rect 8264 36922 8298 37098
rect 8522 36922 8556 37098
rect 8780 36922 8814 37098
rect 9038 36922 9072 37098
rect 9296 36922 9330 37098
rect 9554 36922 9588 37098
rect 9812 36922 9846 37098
rect 10070 36922 10104 37098
rect 10328 36922 10362 37098
rect 10586 36922 10620 37098
rect 12873 36663 12907 36839
rect 13131 36663 13165 36839
rect 13389 36663 13423 36839
rect 20278 37040 20312 37216
rect 20536 37040 20570 37216
rect 20794 37040 20828 37216
rect 21052 37040 21086 37216
rect 21310 37040 21344 37216
rect 21568 37040 21602 37216
rect 21826 37040 21860 37216
rect 22084 37040 22118 37216
rect 22342 37040 22376 37216
rect 22600 37040 22634 37216
rect 22858 37040 22892 37216
rect 23116 37040 23150 37216
rect 23374 37040 23408 37216
rect 12622 35357 12656 35391
rect 12622 35289 12656 35323
rect 12706 35357 12740 35391
rect 12706 35289 12740 35323
rect 12706 35221 12740 35255
rect 12790 35357 12824 35391
rect 12790 35289 12824 35323
rect 12874 35357 12908 35391
rect 12874 35289 12908 35323
rect 12874 35221 12908 35255
rect 12958 35357 12992 35391
rect 12958 35289 12992 35323
rect 13042 35357 13076 35391
rect 13042 35289 13076 35323
rect 13042 35221 13076 35255
rect 13126 35357 13160 35391
rect 13126 35289 13160 35323
rect 13210 35357 13244 35391
rect 13210 35289 13244 35323
rect 13210 35221 13244 35255
rect 13294 35357 13328 35391
rect 13294 35289 13328 35323
rect 25661 36781 25695 36957
rect 25919 36781 25953 36957
rect 26177 36781 26211 36957
rect 25410 35475 25444 35509
rect 25410 35407 25444 35441
rect 25494 35475 25528 35509
rect 25494 35407 25528 35441
rect 25494 35339 25528 35373
rect 25578 35475 25612 35509
rect 25578 35407 25612 35441
rect 25662 35475 25696 35509
rect 25662 35407 25696 35441
rect 25662 35339 25696 35373
rect 25746 35475 25780 35509
rect 25746 35407 25780 35441
rect 25830 35475 25864 35509
rect 25830 35407 25864 35441
rect 25830 35339 25864 35373
rect 25914 35475 25948 35509
rect 25914 35407 25948 35441
rect 25998 35475 26032 35509
rect 25998 35407 26032 35441
rect 25998 35339 26032 35373
rect 26082 35475 26116 35509
rect 26082 35407 26116 35441
rect 12893 32197 12927 32373
rect 13151 32197 13185 32373
rect 13409 32197 13443 32373
rect 25625 32121 25659 32297
rect 25883 32121 25917 32297
rect 26141 32121 26175 32297
rect 7510 30996 7544 31172
rect 7768 30996 7802 31172
rect 8026 30996 8060 31172
rect 8284 30996 8318 31172
rect 8542 30996 8576 31172
rect 8800 30996 8834 31172
rect 9058 30996 9092 31172
rect 9316 30996 9350 31172
rect 9574 30996 9608 31172
rect 9832 30996 9866 31172
rect 10090 30996 10124 31172
rect 10348 30996 10382 31172
rect 10606 30996 10640 31172
rect 12893 30737 12927 30913
rect 13151 30737 13185 30913
rect 13409 30737 13443 30913
rect 12642 29431 12676 29465
rect 12642 29363 12676 29397
rect 12726 29431 12760 29465
rect 12726 29363 12760 29397
rect 12726 29295 12760 29329
rect 12810 29431 12844 29465
rect 12810 29363 12844 29397
rect 12894 29431 12928 29465
rect 12894 29363 12928 29397
rect 12894 29295 12928 29329
rect 12978 29431 13012 29465
rect 12978 29363 13012 29397
rect 13062 29431 13096 29465
rect 13062 29363 13096 29397
rect 13062 29295 13096 29329
rect 13146 29431 13180 29465
rect 13146 29363 13180 29397
rect 13230 29431 13264 29465
rect 13230 29363 13264 29397
rect 13230 29295 13264 29329
rect 13314 29431 13348 29465
rect 13314 29363 13348 29397
rect 20242 30920 20276 31096
rect 20500 30920 20534 31096
rect 20758 30920 20792 31096
rect 21016 30920 21050 31096
rect 21274 30920 21308 31096
rect 21532 30920 21566 31096
rect 21790 30920 21824 31096
rect 22048 30920 22082 31096
rect 22306 30920 22340 31096
rect 22564 30920 22598 31096
rect 22822 30920 22856 31096
rect 23080 30920 23114 31096
rect 23338 30920 23372 31096
rect 25625 30661 25659 30837
rect 25883 30661 25917 30837
rect 26141 30661 26175 30837
rect 25374 29355 25408 29389
rect 25374 29287 25408 29321
rect 25458 29355 25492 29389
rect 25458 29287 25492 29321
rect 25458 29219 25492 29253
rect 25542 29355 25576 29389
rect 25542 29287 25576 29321
rect 25626 29355 25660 29389
rect 25626 29287 25660 29321
rect 25626 29219 25660 29253
rect 25710 29355 25744 29389
rect 25710 29287 25744 29321
rect 25794 29355 25828 29389
rect 25794 29287 25828 29321
rect 25794 29219 25828 29253
rect 25878 29355 25912 29389
rect 25878 29287 25912 29321
rect 25962 29355 25996 29389
rect 25962 29287 25996 29321
rect 25962 29219 25996 29253
rect 26046 29355 26080 29389
rect 26046 29287 26080 29321
rect 13013 25493 13047 25669
rect 13271 25493 13305 25669
rect 13529 25493 13563 25669
rect 25721 25363 25755 25539
rect 25979 25363 26013 25539
rect 26237 25363 26271 25539
rect 7630 24292 7664 24468
rect 7888 24292 7922 24468
rect 8146 24292 8180 24468
rect 8404 24292 8438 24468
rect 8662 24292 8696 24468
rect 8920 24292 8954 24468
rect 9178 24292 9212 24468
rect 9436 24292 9470 24468
rect 9694 24292 9728 24468
rect 9952 24292 9986 24468
rect 10210 24292 10244 24468
rect 10468 24292 10502 24468
rect 10726 24292 10760 24468
rect 13013 24033 13047 24209
rect 13271 24033 13305 24209
rect 13529 24033 13563 24209
rect 12762 22727 12796 22761
rect 12762 22659 12796 22693
rect 12846 22727 12880 22761
rect 12846 22659 12880 22693
rect 12846 22591 12880 22625
rect 12930 22727 12964 22761
rect 12930 22659 12964 22693
rect 13014 22727 13048 22761
rect 13014 22659 13048 22693
rect 13014 22591 13048 22625
rect 13098 22727 13132 22761
rect 13098 22659 13132 22693
rect 13182 22727 13216 22761
rect 13182 22659 13216 22693
rect 13182 22591 13216 22625
rect 13266 22727 13300 22761
rect 13266 22659 13300 22693
rect 13350 22727 13384 22761
rect 13350 22659 13384 22693
rect 13350 22591 13384 22625
rect 13434 22727 13468 22761
rect 13434 22659 13468 22693
rect 20338 24162 20372 24338
rect 20596 24162 20630 24338
rect 20854 24162 20888 24338
rect 21112 24162 21146 24338
rect 21370 24162 21404 24338
rect 21628 24162 21662 24338
rect 21886 24162 21920 24338
rect 22144 24162 22178 24338
rect 22402 24162 22436 24338
rect 22660 24162 22694 24338
rect 22918 24162 22952 24338
rect 23176 24162 23210 24338
rect 23434 24162 23468 24338
rect 25721 23903 25755 24079
rect 25979 23903 26013 24079
rect 26237 23903 26271 24079
rect 25470 22597 25504 22631
rect 25470 22529 25504 22563
rect 25554 22597 25588 22631
rect 25554 22529 25588 22563
rect 25554 22461 25588 22495
rect 25638 22597 25672 22631
rect 25638 22529 25672 22563
rect 25722 22597 25756 22631
rect 25722 22529 25756 22563
rect 25722 22461 25756 22495
rect 25806 22597 25840 22631
rect 25806 22529 25840 22563
rect 25890 22597 25924 22631
rect 25890 22529 25924 22563
rect 25890 22461 25924 22495
rect 25974 22597 26008 22631
rect 25974 22529 26008 22563
rect 26058 22597 26092 22631
rect 26058 22529 26092 22563
rect 26058 22461 26092 22495
rect 26142 22597 26176 22631
rect 26142 22529 26176 22563
rect 12889 18447 12923 18623
rect 13147 18447 13181 18623
rect 13405 18447 13439 18623
rect 26071 18317 26105 18493
rect 26329 18317 26363 18493
rect 26587 18317 26621 18493
rect 7506 17246 7540 17422
rect 7764 17246 7798 17422
rect 8022 17246 8056 17422
rect 8280 17246 8314 17422
rect 8538 17246 8572 17422
rect 8796 17246 8830 17422
rect 9054 17246 9088 17422
rect 9312 17246 9346 17422
rect 9570 17246 9604 17422
rect 9828 17246 9862 17422
rect 10086 17246 10120 17422
rect 10344 17246 10378 17422
rect 10602 17246 10636 17422
rect 12889 16987 12923 17163
rect 13147 16987 13181 17163
rect 13405 16987 13439 17163
rect 12638 15681 12672 15715
rect 12638 15613 12672 15647
rect 12722 15681 12756 15715
rect 12722 15613 12756 15647
rect 12722 15545 12756 15579
rect 12806 15681 12840 15715
rect 12806 15613 12840 15647
rect 12890 15681 12924 15715
rect 12890 15613 12924 15647
rect 12890 15545 12924 15579
rect 12974 15681 13008 15715
rect 12974 15613 13008 15647
rect 13058 15681 13092 15715
rect 13058 15613 13092 15647
rect 13058 15545 13092 15579
rect 13142 15681 13176 15715
rect 13142 15613 13176 15647
rect 13226 15681 13260 15715
rect 13226 15613 13260 15647
rect 13226 15545 13260 15579
rect 13310 15681 13344 15715
rect 13310 15613 13344 15647
rect 20688 17116 20722 17292
rect 20946 17116 20980 17292
rect 21204 17116 21238 17292
rect 21462 17116 21496 17292
rect 21720 17116 21754 17292
rect 21978 17116 22012 17292
rect 22236 17116 22270 17292
rect 22494 17116 22528 17292
rect 22752 17116 22786 17292
rect 23010 17116 23044 17292
rect 23268 17116 23302 17292
rect 23526 17116 23560 17292
rect 23784 17116 23818 17292
rect 26071 16857 26105 17033
rect 26329 16857 26363 17033
rect 26587 16857 26621 17033
rect 25820 15551 25854 15585
rect 25820 15483 25854 15517
rect 25904 15551 25938 15585
rect 25904 15483 25938 15517
rect 25904 15415 25938 15449
rect 25988 15551 26022 15585
rect 25988 15483 26022 15517
rect 26072 15551 26106 15585
rect 26072 15483 26106 15517
rect 26072 15415 26106 15449
rect 26156 15551 26190 15585
rect 26156 15483 26190 15517
rect 26240 15551 26274 15585
rect 26240 15483 26274 15517
rect 26240 15415 26274 15449
rect 26324 15551 26358 15585
rect 26324 15483 26358 15517
rect 26408 15551 26442 15585
rect 26408 15483 26442 15517
rect 26408 15415 26442 15449
rect 26492 15551 26526 15585
rect 26492 15483 26526 15517
<< psubdiff >>
rect 5964 37608 10980 37618
rect 5964 37568 6036 37608
rect 10886 37568 10980 37608
rect 5964 37552 10980 37568
rect 5964 37538 6030 37552
rect 5964 35668 5976 37538
rect 6016 35668 6030 37538
rect 10914 37548 10980 37552
rect 7486 36048 10616 36078
rect 7486 35998 7526 36048
rect 10576 35998 10616 36048
rect 7486 35969 10616 35998
rect 7486 35968 7846 35969
rect 10256 35968 10616 35969
rect 5964 35638 6030 35668
rect 10914 35658 10926 37548
rect 10966 35658 10980 37548
rect 10914 35638 10980 35658
rect 5964 35628 10980 35638
rect 5964 35588 6036 35628
rect 10896 35588 10980 35628
rect 5964 35572 10980 35588
rect 12759 37893 13537 37927
rect 12759 37831 12793 37893
rect 13503 37831 13537 37893
rect 12759 37475 12793 37537
rect 13503 37475 13537 37537
rect 12759 37441 12855 37475
rect 13441 37441 13537 37475
rect 12759 36433 13537 36467
rect 12759 36371 12793 36433
rect 13503 36371 13537 36433
rect 12759 36015 12793 36077
rect 13503 36015 13537 36077
rect 12759 35981 12855 36015
rect 13441 35981 13537 36015
rect 18752 37726 23768 37736
rect 18752 37686 18824 37726
rect 23674 37686 23768 37726
rect 18752 37670 23768 37686
rect 18752 37656 18818 37670
rect 18752 35786 18764 37656
rect 18804 35786 18818 37656
rect 23702 37666 23768 37670
rect 20274 36166 23404 36196
rect 20274 36116 20314 36166
rect 23364 36116 23404 36166
rect 20274 36087 23404 36116
rect 20274 36086 20634 36087
rect 23044 36086 23404 36087
rect 18752 35756 18818 35786
rect 23702 35776 23714 37666
rect 23754 35776 23768 37666
rect 23702 35756 23768 35776
rect 18752 35746 23768 35756
rect 18752 35706 18824 35746
rect 23684 35706 23768 35746
rect 18752 35690 23768 35706
rect 25547 38011 26325 38045
rect 25547 37949 25581 38011
rect 24280 37830 24376 37864
rect 24582 37830 24678 37864
rect 24280 37768 24314 37830
rect 22280 35136 22376 35170
rect 24076 35136 24172 35170
rect 13411 35051 13537 35075
rect 13445 35017 13503 35051
rect 13411 34970 13537 35017
rect 22280 35074 22314 35136
rect 24138 35074 24172 35136
rect 22280 34806 22314 34868
rect 24138 34806 24172 34868
rect 22280 34772 22376 34806
rect 24076 34772 24172 34806
rect 24644 37768 24678 37830
rect 24280 34806 24314 34868
rect 26291 37949 26325 38011
rect 25547 37593 25581 37655
rect 26291 37593 26325 37655
rect 25547 37559 25643 37593
rect 26229 37559 26325 37593
rect 25547 36551 26325 36585
rect 25547 36489 25581 36551
rect 26291 36489 26325 36551
rect 25547 36133 25581 36195
rect 26291 36133 26325 36195
rect 25547 36099 25643 36133
rect 26229 36099 26325 36133
rect 26199 35169 26325 35193
rect 26233 35135 26291 35169
rect 26199 35088 26325 35135
rect 24644 34806 24678 34868
rect 24280 34772 24376 34806
rect 24582 34772 24678 34806
rect 5984 31682 11000 31692
rect 5984 31642 6056 31682
rect 10906 31642 11000 31682
rect 5984 31626 11000 31642
rect 5984 31612 6050 31626
rect 5984 29742 5996 31612
rect 6036 29742 6050 31612
rect 10934 31622 11000 31626
rect 7506 30122 10636 30152
rect 7506 30072 7546 30122
rect 10596 30072 10636 30122
rect 7506 30043 10636 30072
rect 7506 30042 7866 30043
rect 10276 30042 10636 30043
rect 5984 29712 6050 29742
rect 10934 29732 10946 31622
rect 10986 29732 11000 31622
rect 10934 29712 11000 29732
rect 5984 29702 11000 29712
rect 5984 29662 6056 29702
rect 10916 29662 11000 29702
rect 5984 29646 11000 29662
rect 12779 31967 13557 32001
rect 12779 31905 12813 31967
rect 11512 31786 11608 31820
rect 11814 31786 11910 31820
rect 11512 31724 11546 31786
rect 9512 29092 9608 29126
rect 11308 29092 11404 29126
rect 9512 29030 9546 29092
rect 11370 29030 11404 29092
rect 9512 28762 9546 28824
rect 11370 28762 11404 28824
rect 9512 28728 9608 28762
rect 11308 28728 11404 28762
rect 11876 31724 11910 31786
rect 11512 28762 11546 28824
rect 13523 31905 13557 31967
rect 12779 31549 12813 31611
rect 13523 31549 13557 31611
rect 12779 31515 12875 31549
rect 13461 31515 13557 31549
rect 12779 30507 13557 30541
rect 12779 30445 12813 30507
rect 13523 30445 13557 30507
rect 12779 30089 12813 30151
rect 13523 30089 13557 30151
rect 12779 30055 12875 30089
rect 13461 30055 13557 30089
rect 18716 31606 23732 31616
rect 18716 31566 18788 31606
rect 23638 31566 23732 31606
rect 18716 31550 23732 31566
rect 18716 31536 18782 31550
rect 18716 29666 18728 31536
rect 18768 29666 18782 31536
rect 23666 31546 23732 31550
rect 20238 30046 23368 30076
rect 20238 29996 20278 30046
rect 23328 29996 23368 30046
rect 20238 29967 23368 29996
rect 20238 29966 20598 29967
rect 23008 29966 23368 29967
rect 18716 29636 18782 29666
rect 23666 29656 23678 31546
rect 23718 29656 23732 31546
rect 23666 29636 23732 29656
rect 18716 29626 23732 29636
rect 18716 29586 18788 29626
rect 23648 29586 23732 29626
rect 18716 29570 23732 29586
rect 25511 31891 26289 31925
rect 25511 31829 25545 31891
rect 24244 31710 24340 31744
rect 24546 31710 24642 31744
rect 24244 31648 24278 31710
rect 13431 29125 13557 29149
rect 13465 29091 13523 29125
rect 13431 29044 13557 29091
rect 22244 29016 22340 29050
rect 24040 29016 24136 29050
rect 11876 28762 11910 28824
rect 11512 28728 11608 28762
rect 11814 28728 11910 28762
rect 22244 28954 22278 29016
rect 24102 28954 24136 29016
rect 22244 28686 22278 28748
rect 24102 28686 24136 28748
rect 22244 28652 22340 28686
rect 24040 28652 24136 28686
rect 24608 31648 24642 31710
rect 24244 28686 24278 28748
rect 26255 31829 26289 31891
rect 25511 31473 25545 31535
rect 26255 31473 26289 31535
rect 25511 31439 25607 31473
rect 26193 31439 26289 31473
rect 25511 30431 26289 30465
rect 25511 30369 25545 30431
rect 26255 30369 26289 30431
rect 25511 30013 25545 30075
rect 26255 30013 26289 30075
rect 25511 29979 25607 30013
rect 26193 29979 26289 30013
rect 26163 29049 26289 29073
rect 26197 29015 26255 29049
rect 26163 28968 26289 29015
rect 24608 28686 24642 28748
rect 24244 28652 24340 28686
rect 24546 28652 24642 28686
rect 6104 24978 11120 24988
rect 6104 24938 6176 24978
rect 11026 24938 11120 24978
rect 6104 24922 11120 24938
rect 6104 24908 6170 24922
rect 6104 23038 6116 24908
rect 6156 23038 6170 24908
rect 11054 24918 11120 24922
rect 7626 23418 10756 23448
rect 7626 23368 7666 23418
rect 10716 23368 10756 23418
rect 7626 23339 10756 23368
rect 7626 23338 7986 23339
rect 10396 23338 10756 23339
rect 6104 23008 6170 23038
rect 11054 23028 11066 24918
rect 11106 23028 11120 24918
rect 11054 23008 11120 23028
rect 6104 22998 11120 23008
rect 6104 22958 6176 22998
rect 11036 22958 11120 22998
rect 6104 22942 11120 22958
rect 12899 25263 13677 25297
rect 12899 25201 12933 25263
rect 11632 25082 11728 25116
rect 11934 25082 12030 25116
rect 11632 25020 11666 25082
rect 9632 22388 9728 22422
rect 11428 22388 11524 22422
rect 9632 22326 9666 22388
rect 11490 22326 11524 22388
rect 9632 22058 9666 22120
rect 11490 22058 11524 22120
rect 9632 22024 9728 22058
rect 11428 22024 11524 22058
rect 11996 25020 12030 25082
rect 11632 22058 11666 22120
rect 13643 25201 13677 25263
rect 12899 24845 12933 24907
rect 13643 24845 13677 24907
rect 12899 24811 12995 24845
rect 13581 24811 13677 24845
rect 12899 23803 13677 23837
rect 12899 23741 12933 23803
rect 13643 23741 13677 23803
rect 12899 23385 12933 23447
rect 13643 23385 13677 23447
rect 12899 23351 12995 23385
rect 13581 23351 13677 23385
rect 18812 24848 23828 24858
rect 18812 24808 18884 24848
rect 23734 24808 23828 24848
rect 18812 24792 23828 24808
rect 18812 24778 18878 24792
rect 18812 22908 18824 24778
rect 18864 22908 18878 24778
rect 23762 24788 23828 24792
rect 20334 23288 23464 23318
rect 20334 23238 20374 23288
rect 23424 23238 23464 23288
rect 20334 23209 23464 23238
rect 20334 23208 20694 23209
rect 23104 23208 23464 23209
rect 18812 22878 18878 22908
rect 23762 22898 23774 24788
rect 23814 22898 23828 24788
rect 23762 22878 23828 22898
rect 18812 22868 23828 22878
rect 18812 22828 18884 22868
rect 23744 22828 23828 22868
rect 18812 22812 23828 22828
rect 25607 25133 26385 25167
rect 25607 25071 25641 25133
rect 24340 24952 24436 24986
rect 24642 24952 24738 24986
rect 24340 24890 24374 24952
rect 13551 22421 13677 22445
rect 13585 22387 13643 22421
rect 13551 22340 13677 22387
rect 11996 22058 12030 22120
rect 11632 22024 11728 22058
rect 11934 22024 12030 22058
rect 22340 22258 22436 22292
rect 24136 22258 24232 22292
rect 22340 22196 22374 22258
rect 24198 22196 24232 22258
rect 22340 21928 22374 21990
rect 24198 21928 24232 21990
rect 22340 21894 22436 21928
rect 24136 21894 24232 21928
rect 24704 24890 24738 24952
rect 24340 21928 24374 21990
rect 26351 25071 26385 25133
rect 25607 24715 25641 24777
rect 26351 24715 26385 24777
rect 25607 24681 25703 24715
rect 26289 24681 26385 24715
rect 25607 23673 26385 23707
rect 25607 23611 25641 23673
rect 26351 23611 26385 23673
rect 25607 23255 25641 23317
rect 26351 23255 26385 23317
rect 25607 23221 25703 23255
rect 26289 23221 26385 23255
rect 26259 22291 26385 22315
rect 26293 22257 26351 22291
rect 26259 22210 26385 22257
rect 24704 21928 24738 21990
rect 24340 21894 24436 21928
rect 24642 21894 24738 21928
rect 5980 17932 10996 17942
rect 5980 17892 6052 17932
rect 10902 17892 10996 17932
rect 5980 17876 10996 17892
rect 5980 17862 6046 17876
rect 5980 15992 5992 17862
rect 6032 15992 6046 17862
rect 10930 17872 10996 17876
rect 7502 16372 10632 16402
rect 7502 16322 7542 16372
rect 10592 16322 10632 16372
rect 7502 16293 10632 16322
rect 7502 16292 7862 16293
rect 10272 16292 10632 16293
rect 5980 15962 6046 15992
rect 10930 15982 10942 17872
rect 10982 15982 10996 17872
rect 10930 15962 10996 15982
rect 5980 15952 10996 15962
rect 5980 15912 6052 15952
rect 10912 15912 10996 15952
rect 5980 15896 10996 15912
rect 12775 18217 13553 18251
rect 12775 18155 12809 18217
rect 11508 18036 11604 18070
rect 11810 18036 11906 18070
rect 11508 17974 11542 18036
rect 9508 15342 9604 15376
rect 11304 15342 11400 15376
rect 9508 15280 9542 15342
rect 11366 15280 11400 15342
rect 9508 15012 9542 15074
rect 11366 15012 11400 15074
rect 9508 14978 9604 15012
rect 11304 14978 11400 15012
rect 11872 17974 11906 18036
rect 11508 15012 11542 15074
rect 13519 18155 13553 18217
rect 12775 17799 12809 17861
rect 13519 17799 13553 17861
rect 12775 17765 12871 17799
rect 13457 17765 13553 17799
rect 12775 16757 13553 16791
rect 12775 16695 12809 16757
rect 13519 16695 13553 16757
rect 12775 16339 12809 16401
rect 13519 16339 13553 16401
rect 12775 16305 12871 16339
rect 13457 16305 13553 16339
rect 19162 17802 24178 17812
rect 19162 17762 19234 17802
rect 24084 17762 24178 17802
rect 19162 17746 24178 17762
rect 19162 17732 19228 17746
rect 19162 15862 19174 17732
rect 19214 15862 19228 17732
rect 24112 17742 24178 17746
rect 20684 16242 23814 16272
rect 20684 16192 20724 16242
rect 23774 16192 23814 16242
rect 20684 16163 23814 16192
rect 20684 16162 21044 16163
rect 23454 16162 23814 16163
rect 19162 15832 19228 15862
rect 24112 15852 24124 17742
rect 24164 15852 24178 17742
rect 24112 15832 24178 15852
rect 19162 15822 24178 15832
rect 19162 15782 19234 15822
rect 24094 15782 24178 15822
rect 19162 15766 24178 15782
rect 25957 18087 26735 18121
rect 25957 18025 25991 18087
rect 24690 17906 24786 17940
rect 24992 17906 25088 17940
rect 24690 17844 24724 17906
rect 13427 15375 13553 15399
rect 13461 15341 13519 15375
rect 13427 15294 13553 15341
rect 11872 15012 11906 15074
rect 11508 14978 11604 15012
rect 11810 14978 11906 15012
rect 22690 15212 22786 15246
rect 24486 15212 24582 15246
rect 22690 15150 22724 15212
rect 24548 15150 24582 15212
rect 22690 14882 22724 14944
rect 24548 14882 24582 14944
rect 22690 14848 22786 14882
rect 24486 14848 24582 14882
rect 25054 17844 25088 17906
rect 24690 14882 24724 14944
rect 26701 18025 26735 18087
rect 25957 17669 25991 17731
rect 26701 17669 26735 17731
rect 25957 17635 26053 17669
rect 26639 17635 26735 17669
rect 25957 16627 26735 16661
rect 25957 16565 25991 16627
rect 26701 16565 26735 16627
rect 25957 16209 25991 16271
rect 26701 16209 26735 16271
rect 25957 16175 26053 16209
rect 26639 16175 26735 16209
rect 26609 15245 26735 15269
rect 26643 15211 26701 15245
rect 26609 15164 26735 15211
rect 25054 14882 25088 14944
rect 24690 14848 24786 14882
rect 24992 14848 25088 14882
<< nsubdiff >>
rect 25547 38579 25643 38613
rect 26229 38579 26325 38613
rect 25547 38516 25581 38579
rect 12759 38461 12855 38495
rect 13441 38461 13537 38495
rect 12759 38398 12793 38461
rect 13503 38398 13537 38461
rect 12759 38033 12793 38096
rect 26291 38516 26325 38579
rect 25547 38151 25581 38214
rect 26291 38151 26325 38214
rect 25547 38117 26325 38151
rect 13503 38033 13537 38096
rect 12759 37999 13537 38033
rect 18488 38056 24032 38066
rect 18488 38016 18554 38056
rect 23954 38016 24032 38056
rect 18488 38000 24032 38016
rect 18488 37976 18554 38000
rect 5700 37938 11244 37948
rect 5700 37898 5766 37938
rect 11166 37898 11244 37938
rect 5700 37882 11244 37898
rect 5700 37858 5766 37882
rect 5700 35328 5716 37858
rect 5756 35328 5766 37858
rect 11178 37868 11244 37882
rect 7526 37238 10616 37278
rect 7526 37198 7566 37238
rect 10576 37198 10616 37238
rect 7526 37168 10616 37198
rect 5700 35308 5766 35328
rect 11178 35318 11196 37868
rect 11236 35318 11244 37868
rect 12759 37001 12855 37035
rect 13441 37001 13537 37035
rect 12759 36938 12793 37001
rect 13503 36938 13537 37001
rect 12759 36573 12793 36636
rect 13503 36573 13537 36636
rect 12759 36539 13537 36573
rect 18488 35446 18504 37976
rect 18544 35446 18554 37976
rect 23966 37986 24032 38000
rect 20314 37356 23404 37396
rect 20314 37316 20354 37356
rect 23364 37316 23404 37356
rect 20314 37286 23404 37316
rect 18488 35426 18554 35446
rect 23966 35436 23984 37986
rect 24024 35436 24032 37986
rect 23966 35426 24032 35436
rect 18488 35416 24032 35426
rect 11178 35308 11244 35318
rect 5700 35298 11244 35308
rect 5700 35258 5796 35298
rect 11166 35258 11244 35298
rect 5700 35242 11244 35258
rect 13411 35353 13537 35386
rect 18488 35376 18584 35416
rect 23954 35376 24032 35416
rect 18488 35360 24032 35376
rect 13445 35319 13503 35353
rect 13411 35269 13537 35319
rect 13445 35235 13503 35269
rect 13411 35211 13537 35235
rect 25547 37119 25643 37153
rect 26229 37119 26325 37153
rect 25547 37056 25581 37119
rect 26291 37056 26325 37119
rect 25547 36691 25581 36754
rect 26291 36691 26325 36754
rect 25547 36657 26325 36691
rect 26199 35471 26325 35504
rect 26233 35437 26291 35471
rect 26199 35387 26325 35437
rect 26233 35353 26291 35387
rect 26199 35329 26325 35353
rect 12779 32535 12875 32569
rect 13461 32535 13557 32569
rect 12779 32472 12813 32535
rect 13523 32472 13557 32535
rect 12779 32107 12813 32170
rect 13523 32107 13557 32170
rect 12779 32073 13557 32107
rect 25511 32459 25607 32493
rect 26193 32459 26289 32493
rect 25511 32396 25545 32459
rect 26255 32396 26289 32459
rect 25511 32031 25545 32094
rect 26255 32031 26289 32094
rect 5720 32012 11264 32022
rect 5720 31972 5786 32012
rect 11186 31972 11264 32012
rect 5720 31956 11264 31972
rect 5720 31932 5786 31956
rect 5720 29402 5736 31932
rect 5776 29402 5786 31932
rect 11198 31942 11264 31956
rect 7546 31312 10636 31352
rect 7546 31272 7586 31312
rect 10596 31272 10636 31312
rect 7546 31242 10636 31272
rect 5720 29382 5786 29402
rect 11198 29392 11216 31942
rect 11256 29392 11264 31942
rect 25511 31997 26289 32031
rect 11198 29382 11264 29392
rect 5720 29372 11264 29382
rect 5720 29332 5816 29372
rect 11186 29332 11264 29372
rect 5720 29316 11264 29332
rect 18452 31936 23996 31946
rect 18452 31896 18518 31936
rect 23918 31896 23996 31936
rect 18452 31880 23996 31896
rect 18452 31856 18518 31880
rect 12779 31075 12875 31109
rect 13461 31075 13557 31109
rect 12779 31012 12813 31075
rect 13523 31012 13557 31075
rect 12779 30647 12813 30710
rect 13523 30647 13557 30710
rect 12779 30613 13557 30647
rect 13431 29427 13557 29460
rect 13465 29393 13523 29427
rect 13431 29343 13557 29393
rect 13465 29309 13523 29343
rect 13431 29285 13557 29309
rect 18452 29326 18468 31856
rect 18508 29326 18518 31856
rect 23930 31866 23996 31880
rect 20278 31236 23368 31276
rect 20278 31196 20318 31236
rect 23328 31196 23368 31236
rect 20278 31166 23368 31196
rect 18452 29306 18518 29326
rect 23930 29316 23948 31866
rect 23988 29316 23996 31866
rect 23930 29306 23996 29316
rect 18452 29296 23996 29306
rect 18452 29256 18548 29296
rect 23918 29256 23996 29296
rect 18452 29240 23996 29256
rect 25511 30999 25607 31033
rect 26193 30999 26289 31033
rect 25511 30936 25545 30999
rect 26255 30936 26289 30999
rect 25511 30571 25545 30634
rect 26255 30571 26289 30634
rect 25511 30537 26289 30571
rect 26163 29351 26289 29384
rect 26197 29317 26255 29351
rect 26163 29267 26289 29317
rect 26197 29233 26255 29267
rect 26163 29209 26289 29233
rect 12899 25831 12995 25865
rect 13581 25831 13677 25865
rect 12899 25768 12933 25831
rect 13643 25768 13677 25831
rect 12899 25403 12933 25466
rect 13643 25403 13677 25466
rect 12899 25369 13677 25403
rect 25607 25701 25703 25735
rect 26289 25701 26385 25735
rect 25607 25638 25641 25701
rect 26351 25638 26385 25701
rect 5840 25308 11384 25318
rect 5840 25268 5906 25308
rect 11306 25268 11384 25308
rect 5840 25252 11384 25268
rect 5840 25228 5906 25252
rect 5840 22698 5856 25228
rect 5896 22698 5906 25228
rect 11318 25238 11384 25252
rect 7666 24608 10756 24648
rect 7666 24568 7706 24608
rect 10716 24568 10756 24608
rect 7666 24538 10756 24568
rect 5840 22678 5906 22698
rect 11318 22688 11336 25238
rect 11376 22688 11384 25238
rect 11318 22678 11384 22688
rect 5840 22668 11384 22678
rect 5840 22628 5936 22668
rect 11306 22628 11384 22668
rect 5840 22612 11384 22628
rect 25607 25273 25641 25336
rect 26351 25273 26385 25336
rect 25607 25239 26385 25273
rect 18548 25178 24092 25188
rect 18548 25138 18614 25178
rect 24014 25138 24092 25178
rect 18548 25122 24092 25138
rect 18548 25098 18614 25122
rect 12899 24371 12995 24405
rect 13581 24371 13677 24405
rect 12899 24308 12933 24371
rect 13643 24308 13677 24371
rect 12899 23943 12933 24006
rect 13643 23943 13677 24006
rect 12899 23909 13677 23943
rect 13551 22723 13677 22756
rect 13585 22689 13643 22723
rect 13551 22639 13677 22689
rect 13585 22605 13643 22639
rect 13551 22581 13677 22605
rect 18548 22568 18564 25098
rect 18604 22568 18614 25098
rect 24026 25108 24092 25122
rect 20374 24478 23464 24518
rect 20374 24438 20414 24478
rect 23424 24438 23464 24478
rect 20374 24408 23464 24438
rect 18548 22548 18614 22568
rect 24026 22558 24044 25108
rect 24084 22558 24092 25108
rect 24026 22548 24092 22558
rect 18548 22538 24092 22548
rect 18548 22498 18644 22538
rect 24014 22498 24092 22538
rect 18548 22482 24092 22498
rect 25607 24241 25703 24275
rect 26289 24241 26385 24275
rect 25607 24178 25641 24241
rect 26351 24178 26385 24241
rect 25607 23813 25641 23876
rect 26351 23813 26385 23876
rect 25607 23779 26385 23813
rect 26259 22593 26385 22626
rect 26293 22559 26351 22593
rect 26259 22509 26385 22559
rect 26293 22475 26351 22509
rect 26259 22451 26385 22475
rect 12775 18785 12871 18819
rect 13457 18785 13553 18819
rect 12775 18722 12809 18785
rect 13519 18722 13553 18785
rect 12775 18357 12809 18420
rect 13519 18357 13553 18420
rect 12775 18323 13553 18357
rect 25957 18655 26053 18689
rect 26639 18655 26735 18689
rect 25957 18592 25991 18655
rect 26701 18592 26735 18655
rect 5716 18262 11260 18272
rect 5716 18222 5782 18262
rect 11182 18222 11260 18262
rect 5716 18206 11260 18222
rect 5716 18182 5782 18206
rect 5716 15652 5732 18182
rect 5772 15652 5782 18182
rect 11194 18192 11260 18206
rect 7542 17562 10632 17602
rect 7542 17522 7582 17562
rect 10592 17522 10632 17562
rect 7542 17492 10632 17522
rect 5716 15632 5782 15652
rect 11194 15642 11212 18192
rect 11252 15642 11260 18192
rect 11194 15632 11260 15642
rect 5716 15622 11260 15632
rect 5716 15582 5812 15622
rect 11182 15582 11260 15622
rect 5716 15566 11260 15582
rect 25957 18227 25991 18290
rect 26701 18227 26735 18290
rect 25957 18193 26735 18227
rect 18898 18132 24442 18142
rect 18898 18092 18964 18132
rect 24364 18092 24442 18132
rect 18898 18076 24442 18092
rect 18898 18052 18964 18076
rect 12775 17325 12871 17359
rect 13457 17325 13553 17359
rect 12775 17262 12809 17325
rect 13519 17262 13553 17325
rect 12775 16897 12809 16960
rect 13519 16897 13553 16960
rect 12775 16863 13553 16897
rect 13427 15677 13553 15710
rect 13461 15643 13519 15677
rect 13427 15593 13553 15643
rect 13461 15559 13519 15593
rect 13427 15535 13553 15559
rect 18898 15522 18914 18052
rect 18954 15522 18964 18052
rect 24376 18062 24442 18076
rect 20724 17432 23814 17472
rect 20724 17392 20764 17432
rect 23774 17392 23814 17432
rect 20724 17362 23814 17392
rect 18898 15502 18964 15522
rect 24376 15512 24394 18062
rect 24434 15512 24442 18062
rect 24376 15502 24442 15512
rect 18898 15492 24442 15502
rect 18898 15452 18994 15492
rect 24364 15452 24442 15492
rect 18898 15436 24442 15452
rect 25957 17195 26053 17229
rect 26639 17195 26735 17229
rect 25957 17132 25991 17195
rect 26701 17132 26735 17195
rect 25957 16767 25991 16830
rect 26701 16767 26735 16830
rect 25957 16733 26735 16767
rect 26609 15547 26735 15580
rect 26643 15513 26701 15547
rect 26609 15463 26735 15513
rect 26643 15429 26701 15463
rect 26609 15405 26735 15429
<< psubdiffcont >>
rect 6036 37568 10886 37608
rect 5976 35668 6016 37538
rect 7526 35998 10576 36048
rect 10926 35658 10966 37548
rect 6036 35588 10896 35628
rect 12759 37537 12793 37831
rect 13503 37537 13537 37831
rect 12855 37441 13441 37475
rect 12759 36077 12793 36371
rect 13503 36077 13537 36371
rect 12855 35981 13441 36015
rect 18824 37686 23674 37726
rect 18764 35786 18804 37656
rect 20314 36116 23364 36166
rect 23714 35776 23754 37666
rect 18824 35706 23684 35746
rect 24376 37830 24582 37864
rect 22376 35136 24076 35170
rect 13411 35017 13445 35051
rect 13503 35017 13537 35051
rect 22280 34868 22314 35074
rect 24138 34868 24172 35074
rect 22376 34772 24076 34806
rect 24280 34868 24314 37768
rect 24644 34868 24678 37768
rect 25547 37655 25581 37949
rect 26291 37655 26325 37949
rect 25643 37559 26229 37593
rect 25547 36195 25581 36489
rect 26291 36195 26325 36489
rect 25643 36099 26229 36133
rect 26199 35135 26233 35169
rect 26291 35135 26325 35169
rect 24376 34772 24582 34806
rect 6056 31642 10906 31682
rect 5996 29742 6036 31612
rect 7546 30072 10596 30122
rect 10946 29732 10986 31622
rect 6056 29662 10916 29702
rect 11608 31786 11814 31820
rect 9608 29092 11308 29126
rect 9512 28824 9546 29030
rect 11370 28824 11404 29030
rect 9608 28728 11308 28762
rect 11512 28824 11546 31724
rect 11876 28824 11910 31724
rect 12779 31611 12813 31905
rect 13523 31611 13557 31905
rect 12875 31515 13461 31549
rect 12779 30151 12813 30445
rect 13523 30151 13557 30445
rect 12875 30055 13461 30089
rect 18788 31566 23638 31606
rect 18728 29666 18768 31536
rect 20278 29996 23328 30046
rect 23678 29656 23718 31546
rect 18788 29586 23648 29626
rect 24340 31710 24546 31744
rect 13431 29091 13465 29125
rect 13523 29091 13557 29125
rect 22340 29016 24040 29050
rect 11608 28728 11814 28762
rect 22244 28748 22278 28954
rect 24102 28748 24136 28954
rect 22340 28652 24040 28686
rect 24244 28748 24278 31648
rect 24608 28748 24642 31648
rect 25511 31535 25545 31829
rect 26255 31535 26289 31829
rect 25607 31439 26193 31473
rect 25511 30075 25545 30369
rect 26255 30075 26289 30369
rect 25607 29979 26193 30013
rect 26163 29015 26197 29049
rect 26255 29015 26289 29049
rect 24340 28652 24546 28686
rect 6176 24938 11026 24978
rect 6116 23038 6156 24908
rect 7666 23368 10716 23418
rect 11066 23028 11106 24918
rect 6176 22958 11036 22998
rect 11728 25082 11934 25116
rect 9728 22388 11428 22422
rect 9632 22120 9666 22326
rect 11490 22120 11524 22326
rect 9728 22024 11428 22058
rect 11632 22120 11666 25020
rect 11996 22120 12030 25020
rect 12899 24907 12933 25201
rect 13643 24907 13677 25201
rect 12995 24811 13581 24845
rect 12899 23447 12933 23741
rect 13643 23447 13677 23741
rect 12995 23351 13581 23385
rect 18884 24808 23734 24848
rect 18824 22908 18864 24778
rect 20374 23238 23424 23288
rect 23774 22898 23814 24788
rect 18884 22828 23744 22868
rect 24436 24952 24642 24986
rect 13551 22387 13585 22421
rect 13643 22387 13677 22421
rect 11728 22024 11934 22058
rect 22436 22258 24136 22292
rect 22340 21990 22374 22196
rect 24198 21990 24232 22196
rect 22436 21894 24136 21928
rect 24340 21990 24374 24890
rect 24704 21990 24738 24890
rect 25607 24777 25641 25071
rect 26351 24777 26385 25071
rect 25703 24681 26289 24715
rect 25607 23317 25641 23611
rect 26351 23317 26385 23611
rect 25703 23221 26289 23255
rect 26259 22257 26293 22291
rect 26351 22257 26385 22291
rect 24436 21894 24642 21928
rect 6052 17892 10902 17932
rect 5992 15992 6032 17862
rect 7542 16322 10592 16372
rect 10942 15982 10982 17872
rect 6052 15912 10912 15952
rect 11604 18036 11810 18070
rect 9604 15342 11304 15376
rect 9508 15074 9542 15280
rect 11366 15074 11400 15280
rect 9604 14978 11304 15012
rect 11508 15074 11542 17974
rect 11872 15074 11906 17974
rect 12775 17861 12809 18155
rect 13519 17861 13553 18155
rect 12871 17765 13457 17799
rect 12775 16401 12809 16695
rect 13519 16401 13553 16695
rect 12871 16305 13457 16339
rect 19234 17762 24084 17802
rect 19174 15862 19214 17732
rect 20724 16192 23774 16242
rect 24124 15852 24164 17742
rect 19234 15782 24094 15822
rect 24786 17906 24992 17940
rect 13427 15341 13461 15375
rect 13519 15341 13553 15375
rect 11604 14978 11810 15012
rect 22786 15212 24486 15246
rect 22690 14944 22724 15150
rect 24548 14944 24582 15150
rect 22786 14848 24486 14882
rect 24690 14944 24724 17844
rect 25054 14944 25088 17844
rect 25957 17731 25991 18025
rect 26701 17731 26735 18025
rect 26053 17635 26639 17669
rect 25957 16271 25991 16565
rect 26701 16271 26735 16565
rect 26053 16175 26639 16209
rect 26609 15211 26643 15245
rect 26701 15211 26735 15245
rect 24786 14848 24992 14882
<< nsubdiffcont >>
rect 25643 38579 26229 38613
rect 12855 38461 13441 38495
rect 12759 38096 12793 38398
rect 13503 38096 13537 38398
rect 25547 38214 25581 38516
rect 26291 38214 26325 38516
rect 18554 38016 23954 38056
rect 5766 37898 11166 37938
rect 5716 35328 5756 37858
rect 7566 37198 10576 37238
rect 11196 35318 11236 37868
rect 12855 37001 13441 37035
rect 12759 36636 12793 36938
rect 13503 36636 13537 36938
rect 18504 35446 18544 37976
rect 20354 37316 23364 37356
rect 23984 35436 24024 37986
rect 5796 35258 11166 35298
rect 18584 35376 23954 35416
rect 13411 35319 13445 35353
rect 13503 35319 13537 35353
rect 13411 35235 13445 35269
rect 13503 35235 13537 35269
rect 25643 37119 26229 37153
rect 25547 36754 25581 37056
rect 26291 36754 26325 37056
rect 26199 35437 26233 35471
rect 26291 35437 26325 35471
rect 26199 35353 26233 35387
rect 26291 35353 26325 35387
rect 12875 32535 13461 32569
rect 12779 32170 12813 32472
rect 13523 32170 13557 32472
rect 25607 32459 26193 32493
rect 25511 32094 25545 32396
rect 26255 32094 26289 32396
rect 5786 31972 11186 32012
rect 5736 29402 5776 31932
rect 7586 31272 10596 31312
rect 11216 29392 11256 31942
rect 5816 29332 11186 29372
rect 18518 31896 23918 31936
rect 12875 31075 13461 31109
rect 12779 30710 12813 31012
rect 13523 30710 13557 31012
rect 13431 29393 13465 29427
rect 13523 29393 13557 29427
rect 13431 29309 13465 29343
rect 13523 29309 13557 29343
rect 18468 29326 18508 31856
rect 20318 31196 23328 31236
rect 23948 29316 23988 31866
rect 18548 29256 23918 29296
rect 25607 30999 26193 31033
rect 25511 30634 25545 30936
rect 26255 30634 26289 30936
rect 26163 29317 26197 29351
rect 26255 29317 26289 29351
rect 26163 29233 26197 29267
rect 26255 29233 26289 29267
rect 12995 25831 13581 25865
rect 12899 25466 12933 25768
rect 13643 25466 13677 25768
rect 25703 25701 26289 25735
rect 25607 25336 25641 25638
rect 5906 25268 11306 25308
rect 5856 22698 5896 25228
rect 7706 24568 10716 24608
rect 11336 22688 11376 25238
rect 5936 22628 11306 22668
rect 26351 25336 26385 25638
rect 18614 25138 24014 25178
rect 12995 24371 13581 24405
rect 12899 24006 12933 24308
rect 13643 24006 13677 24308
rect 13551 22689 13585 22723
rect 13643 22689 13677 22723
rect 13551 22605 13585 22639
rect 13643 22605 13677 22639
rect 18564 22568 18604 25098
rect 20414 24438 23424 24478
rect 24044 22558 24084 25108
rect 18644 22498 24014 22538
rect 25703 24241 26289 24275
rect 25607 23876 25641 24178
rect 26351 23876 26385 24178
rect 26259 22559 26293 22593
rect 26351 22559 26385 22593
rect 26259 22475 26293 22509
rect 26351 22475 26385 22509
rect 12871 18785 13457 18819
rect 12775 18420 12809 18722
rect 13519 18420 13553 18722
rect 26053 18655 26639 18689
rect 25957 18290 25991 18592
rect 5782 18222 11182 18262
rect 5732 15652 5772 18182
rect 7582 17522 10592 17562
rect 11212 15642 11252 18192
rect 5812 15582 11182 15622
rect 26701 18290 26735 18592
rect 18964 18092 24364 18132
rect 12871 17325 13457 17359
rect 12775 16960 12809 17262
rect 13519 16960 13553 17262
rect 13427 15643 13461 15677
rect 13519 15643 13553 15677
rect 13427 15559 13461 15593
rect 13519 15559 13553 15593
rect 18914 15522 18954 18052
rect 20764 17392 23774 17432
rect 24394 15512 24434 18062
rect 18994 15452 24364 15492
rect 26053 17195 26639 17229
rect 25957 16830 25991 17132
rect 26701 16830 26735 17132
rect 26609 15513 26643 15547
rect 26701 15513 26735 15547
rect 26609 15429 26643 15463
rect 26701 15429 26735 15463
<< poly >>
rect 12919 38392 13119 38408
rect 12919 38358 12935 38392
rect 13103 38358 13119 38392
rect 12919 38311 13119 38358
rect 13177 38392 13377 38408
rect 13177 38358 13193 38392
rect 13361 38358 13377 38392
rect 13177 38311 13377 38358
rect 12919 38085 13119 38111
rect 13177 38085 13377 38111
rect 25707 38510 25907 38526
rect 25707 38476 25723 38510
rect 25891 38476 25907 38510
rect 25707 38429 25907 38476
rect 25965 38510 26165 38526
rect 25965 38476 25981 38510
rect 26149 38476 26165 38510
rect 25965 38429 26165 38476
rect 25707 38203 25907 38229
rect 25965 38203 26165 38229
rect 7536 37110 7736 37136
rect 7794 37110 7994 37136
rect 8052 37110 8252 37136
rect 8310 37110 8510 37136
rect 8568 37110 8768 37136
rect 8826 37110 9026 37136
rect 9084 37110 9284 37136
rect 9342 37110 9542 37136
rect 9600 37110 9800 37136
rect 9858 37110 10058 37136
rect 10116 37110 10316 37136
rect 10374 37110 10574 37136
rect 7536 36863 7736 36910
rect 7536 36829 7552 36863
rect 7720 36829 7736 36863
rect 7536 36813 7736 36829
rect 7794 36863 7994 36910
rect 7794 36829 7810 36863
rect 7978 36829 7994 36863
rect 7794 36813 7994 36829
rect 8052 36863 8252 36910
rect 8052 36829 8068 36863
rect 8236 36829 8252 36863
rect 8052 36813 8252 36829
rect 8310 36863 8510 36910
rect 8310 36829 8326 36863
rect 8494 36829 8510 36863
rect 8310 36813 8510 36829
rect 8568 36863 8768 36910
rect 8568 36829 8584 36863
rect 8752 36829 8768 36863
rect 8568 36813 8768 36829
rect 8826 36863 9026 36910
rect 8826 36829 8842 36863
rect 9010 36829 9026 36863
rect 8826 36813 9026 36829
rect 9084 36863 9284 36910
rect 9084 36829 9100 36863
rect 9268 36829 9284 36863
rect 9084 36813 9284 36829
rect 9342 36863 9542 36910
rect 9342 36829 9358 36863
rect 9526 36829 9542 36863
rect 9342 36813 9542 36829
rect 9600 36863 9800 36910
rect 9600 36829 9616 36863
rect 9784 36829 9800 36863
rect 9600 36813 9800 36829
rect 9858 36863 10058 36910
rect 9858 36829 9874 36863
rect 10042 36829 10058 36863
rect 9858 36813 10058 36829
rect 10116 36863 10316 36910
rect 10116 36829 10132 36863
rect 10300 36829 10316 36863
rect 10116 36813 10316 36829
rect 10374 36863 10574 36910
rect 10374 36829 10390 36863
rect 10558 36829 10574 36863
rect 10374 36813 10574 36829
rect 7794 36755 7994 36771
rect 7794 36721 7810 36755
rect 7978 36721 7994 36755
rect 7536 36683 7736 36709
rect 7794 36683 7994 36721
rect 8568 36755 8768 36771
rect 8568 36721 8584 36755
rect 8752 36721 8768 36755
rect 8052 36683 8252 36709
rect 8310 36683 8510 36709
rect 8568 36683 8768 36721
rect 8826 36755 9026 36771
rect 8826 36721 8842 36755
rect 9010 36721 9026 36755
rect 8826 36683 9026 36721
rect 9600 36755 9800 36771
rect 9600 36721 9616 36755
rect 9784 36721 9800 36755
rect 9084 36683 9284 36709
rect 9342 36683 9542 36709
rect 9600 36683 9800 36721
rect 9858 36755 10058 36771
rect 9858 36721 9874 36755
rect 10042 36721 10058 36755
rect 9858 36683 10058 36721
rect 10116 36683 10316 36709
rect 10374 36683 10574 36709
rect 7536 36445 7736 36483
rect 7794 36457 7994 36483
rect 7536 36411 7552 36445
rect 7720 36411 7736 36445
rect 7536 36395 7736 36411
rect 8052 36445 8252 36483
rect 8052 36411 8068 36445
rect 8236 36411 8252 36445
rect 8052 36395 8252 36411
rect 8310 36445 8510 36483
rect 8568 36457 8768 36483
rect 8826 36457 9026 36483
rect 8310 36411 8326 36445
rect 8494 36411 8510 36445
rect 8310 36395 8510 36411
rect 9084 36445 9284 36483
rect 9084 36411 9100 36445
rect 9268 36411 9284 36445
rect 9084 36395 9284 36411
rect 9342 36445 9542 36483
rect 9600 36457 9800 36483
rect 9858 36457 10058 36483
rect 9342 36411 9358 36445
rect 9526 36411 9542 36445
rect 9342 36395 9542 36411
rect 10116 36445 10316 36483
rect 10116 36411 10132 36445
rect 10300 36411 10316 36445
rect 10116 36395 10316 36411
rect 10374 36445 10574 36483
rect 10374 36411 10390 36445
rect 10558 36411 10574 36445
rect 10374 36395 10574 36411
rect 7536 36319 7736 36335
rect 7536 36285 7552 36319
rect 7720 36285 7736 36319
rect 7536 36247 7736 36285
rect 7794 36319 7994 36335
rect 7794 36285 7810 36319
rect 7978 36285 7994 36319
rect 7794 36247 7994 36285
rect 8052 36319 8252 36335
rect 8052 36285 8068 36319
rect 8236 36285 8252 36319
rect 8052 36247 8252 36285
rect 8310 36319 8510 36335
rect 8310 36285 8326 36319
rect 8494 36285 8510 36319
rect 8310 36247 8510 36285
rect 8568 36319 8768 36335
rect 8568 36285 8584 36319
rect 8752 36285 8768 36319
rect 8568 36247 8768 36285
rect 8826 36319 9026 36335
rect 8826 36285 8842 36319
rect 9010 36285 9026 36319
rect 8826 36247 9026 36285
rect 9084 36319 9284 36335
rect 9084 36285 9100 36319
rect 9268 36285 9284 36319
rect 9084 36247 9284 36285
rect 9342 36319 9542 36335
rect 9342 36285 9358 36319
rect 9526 36285 9542 36319
rect 9342 36247 9542 36285
rect 9600 36319 9800 36335
rect 9600 36285 9616 36319
rect 9784 36285 9800 36319
rect 9600 36247 9800 36285
rect 9858 36319 10058 36335
rect 9858 36285 9874 36319
rect 10042 36285 10058 36319
rect 9858 36247 10058 36285
rect 10116 36319 10316 36335
rect 10116 36285 10132 36319
rect 10300 36285 10316 36319
rect 10116 36247 10316 36285
rect 10374 36319 10574 36335
rect 10374 36285 10390 36319
rect 10558 36285 10574 36319
rect 10374 36247 10574 36285
rect 7536 36137 7736 36163
rect 7794 36137 7994 36163
rect 8052 36137 8252 36163
rect 8310 36137 8510 36163
rect 8568 36137 8768 36163
rect 8826 36137 9026 36163
rect 9084 36137 9284 36163
rect 9342 36137 9542 36163
rect 9600 36137 9800 36163
rect 9858 36137 10058 36163
rect 10116 36137 10316 36163
rect 10374 36137 10574 36163
rect 12919 37815 13119 37841
rect 13177 37815 13377 37841
rect 12919 37577 13119 37615
rect 12919 37543 12935 37577
rect 13103 37543 13119 37577
rect 12919 37527 13119 37543
rect 13177 37577 13377 37615
rect 13177 37543 13193 37577
rect 13361 37543 13377 37577
rect 13177 37527 13377 37543
rect 12919 36932 13119 36948
rect 12919 36898 12935 36932
rect 13103 36898 13119 36932
rect 12919 36851 13119 36898
rect 13177 36932 13377 36948
rect 13177 36898 13193 36932
rect 13361 36898 13377 36932
rect 13177 36851 13377 36898
rect 12919 36625 13119 36651
rect 13177 36625 13377 36651
rect 12919 36355 13119 36381
rect 13177 36355 13377 36381
rect 12919 36117 13119 36155
rect 12919 36083 12935 36117
rect 13103 36083 13119 36117
rect 12919 36067 13119 36083
rect 13177 36117 13377 36155
rect 13177 36083 13193 36117
rect 13361 36083 13377 36117
rect 13177 36067 13377 36083
rect 20324 37228 20524 37254
rect 20582 37228 20782 37254
rect 20840 37228 21040 37254
rect 21098 37228 21298 37254
rect 21356 37228 21556 37254
rect 21614 37228 21814 37254
rect 21872 37228 22072 37254
rect 22130 37228 22330 37254
rect 22388 37228 22588 37254
rect 22646 37228 22846 37254
rect 22904 37228 23104 37254
rect 23162 37228 23362 37254
rect 20324 36981 20524 37028
rect 20324 36947 20340 36981
rect 20508 36947 20524 36981
rect 20324 36931 20524 36947
rect 20582 36981 20782 37028
rect 20582 36947 20598 36981
rect 20766 36947 20782 36981
rect 20582 36931 20782 36947
rect 20840 36981 21040 37028
rect 20840 36947 20856 36981
rect 21024 36947 21040 36981
rect 20840 36931 21040 36947
rect 21098 36981 21298 37028
rect 21098 36947 21114 36981
rect 21282 36947 21298 36981
rect 21098 36931 21298 36947
rect 21356 36981 21556 37028
rect 21356 36947 21372 36981
rect 21540 36947 21556 36981
rect 21356 36931 21556 36947
rect 21614 36981 21814 37028
rect 21614 36947 21630 36981
rect 21798 36947 21814 36981
rect 21614 36931 21814 36947
rect 21872 36981 22072 37028
rect 21872 36947 21888 36981
rect 22056 36947 22072 36981
rect 21872 36931 22072 36947
rect 22130 36981 22330 37028
rect 22130 36947 22146 36981
rect 22314 36947 22330 36981
rect 22130 36931 22330 36947
rect 22388 36981 22588 37028
rect 22388 36947 22404 36981
rect 22572 36947 22588 36981
rect 22388 36931 22588 36947
rect 22646 36981 22846 37028
rect 22646 36947 22662 36981
rect 22830 36947 22846 36981
rect 22646 36931 22846 36947
rect 22904 36981 23104 37028
rect 22904 36947 22920 36981
rect 23088 36947 23104 36981
rect 22904 36931 23104 36947
rect 23162 36981 23362 37028
rect 23162 36947 23178 36981
rect 23346 36947 23362 36981
rect 23162 36931 23362 36947
rect 20582 36873 20782 36889
rect 20582 36839 20598 36873
rect 20766 36839 20782 36873
rect 20324 36801 20524 36827
rect 20582 36801 20782 36839
rect 21356 36873 21556 36889
rect 21356 36839 21372 36873
rect 21540 36839 21556 36873
rect 20840 36801 21040 36827
rect 21098 36801 21298 36827
rect 21356 36801 21556 36839
rect 21614 36873 21814 36889
rect 21614 36839 21630 36873
rect 21798 36839 21814 36873
rect 21614 36801 21814 36839
rect 22388 36873 22588 36889
rect 22388 36839 22404 36873
rect 22572 36839 22588 36873
rect 21872 36801 22072 36827
rect 22130 36801 22330 36827
rect 22388 36801 22588 36839
rect 22646 36873 22846 36889
rect 22646 36839 22662 36873
rect 22830 36839 22846 36873
rect 22646 36801 22846 36839
rect 22904 36801 23104 36827
rect 23162 36801 23362 36827
rect 20324 36563 20524 36601
rect 20582 36575 20782 36601
rect 20324 36529 20340 36563
rect 20508 36529 20524 36563
rect 20324 36513 20524 36529
rect 20840 36563 21040 36601
rect 20840 36529 20856 36563
rect 21024 36529 21040 36563
rect 20840 36513 21040 36529
rect 21098 36563 21298 36601
rect 21356 36575 21556 36601
rect 21614 36575 21814 36601
rect 21098 36529 21114 36563
rect 21282 36529 21298 36563
rect 21098 36513 21298 36529
rect 21872 36563 22072 36601
rect 21872 36529 21888 36563
rect 22056 36529 22072 36563
rect 21872 36513 22072 36529
rect 22130 36563 22330 36601
rect 22388 36575 22588 36601
rect 22646 36575 22846 36601
rect 22130 36529 22146 36563
rect 22314 36529 22330 36563
rect 22130 36513 22330 36529
rect 22904 36563 23104 36601
rect 22904 36529 22920 36563
rect 23088 36529 23104 36563
rect 22904 36513 23104 36529
rect 23162 36563 23362 36601
rect 23162 36529 23178 36563
rect 23346 36529 23362 36563
rect 23162 36513 23362 36529
rect 20324 36437 20524 36453
rect 20324 36403 20340 36437
rect 20508 36403 20524 36437
rect 20324 36365 20524 36403
rect 20582 36437 20782 36453
rect 20582 36403 20598 36437
rect 20766 36403 20782 36437
rect 20582 36365 20782 36403
rect 20840 36437 21040 36453
rect 20840 36403 20856 36437
rect 21024 36403 21040 36437
rect 20840 36365 21040 36403
rect 21098 36437 21298 36453
rect 21098 36403 21114 36437
rect 21282 36403 21298 36437
rect 21098 36365 21298 36403
rect 21356 36437 21556 36453
rect 21356 36403 21372 36437
rect 21540 36403 21556 36437
rect 21356 36365 21556 36403
rect 21614 36437 21814 36453
rect 21614 36403 21630 36437
rect 21798 36403 21814 36437
rect 21614 36365 21814 36403
rect 21872 36437 22072 36453
rect 21872 36403 21888 36437
rect 22056 36403 22072 36437
rect 21872 36365 22072 36403
rect 22130 36437 22330 36453
rect 22130 36403 22146 36437
rect 22314 36403 22330 36437
rect 22130 36365 22330 36403
rect 22388 36437 22588 36453
rect 22388 36403 22404 36437
rect 22572 36403 22588 36437
rect 22388 36365 22588 36403
rect 22646 36437 22846 36453
rect 22646 36403 22662 36437
rect 22830 36403 22846 36437
rect 22646 36365 22846 36403
rect 22904 36437 23104 36453
rect 22904 36403 22920 36437
rect 23088 36403 23104 36437
rect 22904 36365 23104 36403
rect 23162 36437 23362 36453
rect 23162 36403 23178 36437
rect 23346 36403 23362 36437
rect 23162 36365 23362 36403
rect 20324 36255 20524 36281
rect 20582 36255 20782 36281
rect 20840 36255 21040 36281
rect 21098 36255 21298 36281
rect 21356 36255 21556 36281
rect 21614 36255 21814 36281
rect 21872 36255 22072 36281
rect 22130 36255 22330 36281
rect 22388 36255 22588 36281
rect 22646 36255 22846 36281
rect 22904 36255 23104 36281
rect 23162 36255 23362 36281
rect 12666 35403 12696 35429
rect 12750 35403 12780 35429
rect 12834 35403 12864 35429
rect 12918 35403 12948 35429
rect 13002 35403 13032 35429
rect 13086 35403 13116 35429
rect 13170 35403 13200 35429
rect 13254 35403 13284 35429
rect 12666 35171 12696 35203
rect 12750 35171 12780 35203
rect 12834 35171 12864 35203
rect 12918 35171 12948 35203
rect 13002 35171 13032 35203
rect 13086 35171 13116 35203
rect 13170 35171 13200 35203
rect 13254 35171 13284 35203
rect 12666 35155 13284 35171
rect 12666 35121 12706 35155
rect 12740 35121 12790 35155
rect 12824 35121 12874 35155
rect 12908 35121 12958 35155
rect 12992 35121 13042 35155
rect 13076 35121 13126 35155
rect 13160 35121 13210 35155
rect 13244 35121 13284 35155
rect 12666 35105 13284 35121
rect 12666 35083 12696 35105
rect 12750 35083 12780 35105
rect 12834 35083 12864 35105
rect 12918 35083 12948 35105
rect 13002 35083 13032 35105
rect 13086 35083 13116 35105
rect 13170 35083 13200 35105
rect 13254 35083 13284 35105
rect 12666 34927 12696 34953
rect 12750 34927 12780 34953
rect 12834 34927 12864 34953
rect 12918 34927 12948 34953
rect 13002 34927 13032 34953
rect 13086 34927 13116 34953
rect 13170 34927 13200 34953
rect 13254 34927 13284 34953
rect 25707 37933 25907 37959
rect 25965 37933 26165 37959
rect 25707 37695 25907 37733
rect 25707 37661 25723 37695
rect 25891 37661 25907 37695
rect 25707 37645 25907 37661
rect 25965 37695 26165 37733
rect 25965 37661 25981 37695
rect 26149 37661 26165 37695
rect 25965 37645 26165 37661
rect 25707 37050 25907 37066
rect 25707 37016 25723 37050
rect 25891 37016 25907 37050
rect 25707 36969 25907 37016
rect 25965 37050 26165 37066
rect 25965 37016 25981 37050
rect 26149 37016 26165 37050
rect 25965 36969 26165 37016
rect 25707 36743 25907 36769
rect 25965 36743 26165 36769
rect 25707 36473 25907 36499
rect 25965 36473 26165 36499
rect 25707 36235 25907 36273
rect 25707 36201 25723 36235
rect 25891 36201 25907 36235
rect 25707 36185 25907 36201
rect 25965 36235 26165 36273
rect 25965 36201 25981 36235
rect 26149 36201 26165 36235
rect 25965 36185 26165 36201
rect 25454 35521 25484 35547
rect 25538 35521 25568 35547
rect 25622 35521 25652 35547
rect 25706 35521 25736 35547
rect 25790 35521 25820 35547
rect 25874 35521 25904 35547
rect 25958 35521 25988 35547
rect 26042 35521 26072 35547
rect 25454 35289 25484 35321
rect 25538 35289 25568 35321
rect 25622 35289 25652 35321
rect 25706 35289 25736 35321
rect 25790 35289 25820 35321
rect 25874 35289 25904 35321
rect 25958 35289 25988 35321
rect 26042 35289 26072 35321
rect 25454 35273 26072 35289
rect 25454 35239 25494 35273
rect 25528 35239 25578 35273
rect 25612 35239 25662 35273
rect 25696 35239 25746 35273
rect 25780 35239 25830 35273
rect 25864 35239 25914 35273
rect 25948 35239 25998 35273
rect 26032 35239 26072 35273
rect 25454 35223 26072 35239
rect 25454 35201 25484 35223
rect 25538 35201 25568 35223
rect 25622 35201 25652 35223
rect 25706 35201 25736 35223
rect 25790 35201 25820 35223
rect 25874 35201 25904 35223
rect 25958 35201 25988 35223
rect 26042 35201 26072 35223
rect 25454 35045 25484 35071
rect 25538 35045 25568 35071
rect 25622 35045 25652 35071
rect 25706 35045 25736 35071
rect 25790 35045 25820 35071
rect 25874 35045 25904 35071
rect 25958 35045 25988 35071
rect 26042 35045 26072 35071
rect 12939 32466 13139 32482
rect 12939 32432 12955 32466
rect 13123 32432 13139 32466
rect 12939 32385 13139 32432
rect 13197 32466 13397 32482
rect 13197 32432 13213 32466
rect 13381 32432 13397 32466
rect 13197 32385 13397 32432
rect 12939 32159 13139 32185
rect 13197 32159 13397 32185
rect 25671 32390 25871 32406
rect 25671 32356 25687 32390
rect 25855 32356 25871 32390
rect 25671 32309 25871 32356
rect 25929 32390 26129 32406
rect 25929 32356 25945 32390
rect 26113 32356 26129 32390
rect 25929 32309 26129 32356
rect 25671 32083 25871 32109
rect 25929 32083 26129 32109
rect 7556 31184 7756 31210
rect 7814 31184 8014 31210
rect 8072 31184 8272 31210
rect 8330 31184 8530 31210
rect 8588 31184 8788 31210
rect 8846 31184 9046 31210
rect 9104 31184 9304 31210
rect 9362 31184 9562 31210
rect 9620 31184 9820 31210
rect 9878 31184 10078 31210
rect 10136 31184 10336 31210
rect 10394 31184 10594 31210
rect 7556 30937 7756 30984
rect 7556 30903 7572 30937
rect 7740 30903 7756 30937
rect 7556 30887 7756 30903
rect 7814 30937 8014 30984
rect 7814 30903 7830 30937
rect 7998 30903 8014 30937
rect 7814 30887 8014 30903
rect 8072 30937 8272 30984
rect 8072 30903 8088 30937
rect 8256 30903 8272 30937
rect 8072 30887 8272 30903
rect 8330 30937 8530 30984
rect 8330 30903 8346 30937
rect 8514 30903 8530 30937
rect 8330 30887 8530 30903
rect 8588 30937 8788 30984
rect 8588 30903 8604 30937
rect 8772 30903 8788 30937
rect 8588 30887 8788 30903
rect 8846 30937 9046 30984
rect 8846 30903 8862 30937
rect 9030 30903 9046 30937
rect 8846 30887 9046 30903
rect 9104 30937 9304 30984
rect 9104 30903 9120 30937
rect 9288 30903 9304 30937
rect 9104 30887 9304 30903
rect 9362 30937 9562 30984
rect 9362 30903 9378 30937
rect 9546 30903 9562 30937
rect 9362 30887 9562 30903
rect 9620 30937 9820 30984
rect 9620 30903 9636 30937
rect 9804 30903 9820 30937
rect 9620 30887 9820 30903
rect 9878 30937 10078 30984
rect 9878 30903 9894 30937
rect 10062 30903 10078 30937
rect 9878 30887 10078 30903
rect 10136 30937 10336 30984
rect 10136 30903 10152 30937
rect 10320 30903 10336 30937
rect 10136 30887 10336 30903
rect 10394 30937 10594 30984
rect 10394 30903 10410 30937
rect 10578 30903 10594 30937
rect 10394 30887 10594 30903
rect 7814 30829 8014 30845
rect 7814 30795 7830 30829
rect 7998 30795 8014 30829
rect 7556 30757 7756 30783
rect 7814 30757 8014 30795
rect 8588 30829 8788 30845
rect 8588 30795 8604 30829
rect 8772 30795 8788 30829
rect 8072 30757 8272 30783
rect 8330 30757 8530 30783
rect 8588 30757 8788 30795
rect 8846 30829 9046 30845
rect 8846 30795 8862 30829
rect 9030 30795 9046 30829
rect 8846 30757 9046 30795
rect 9620 30829 9820 30845
rect 9620 30795 9636 30829
rect 9804 30795 9820 30829
rect 9104 30757 9304 30783
rect 9362 30757 9562 30783
rect 9620 30757 9820 30795
rect 9878 30829 10078 30845
rect 9878 30795 9894 30829
rect 10062 30795 10078 30829
rect 9878 30757 10078 30795
rect 10136 30757 10336 30783
rect 10394 30757 10594 30783
rect 7556 30519 7756 30557
rect 7814 30531 8014 30557
rect 7556 30485 7572 30519
rect 7740 30485 7756 30519
rect 7556 30469 7756 30485
rect 8072 30519 8272 30557
rect 8072 30485 8088 30519
rect 8256 30485 8272 30519
rect 8072 30469 8272 30485
rect 8330 30519 8530 30557
rect 8588 30531 8788 30557
rect 8846 30531 9046 30557
rect 8330 30485 8346 30519
rect 8514 30485 8530 30519
rect 8330 30469 8530 30485
rect 9104 30519 9304 30557
rect 9104 30485 9120 30519
rect 9288 30485 9304 30519
rect 9104 30469 9304 30485
rect 9362 30519 9562 30557
rect 9620 30531 9820 30557
rect 9878 30531 10078 30557
rect 9362 30485 9378 30519
rect 9546 30485 9562 30519
rect 9362 30469 9562 30485
rect 10136 30519 10336 30557
rect 10136 30485 10152 30519
rect 10320 30485 10336 30519
rect 10136 30469 10336 30485
rect 10394 30519 10594 30557
rect 10394 30485 10410 30519
rect 10578 30485 10594 30519
rect 10394 30469 10594 30485
rect 7556 30393 7756 30409
rect 7556 30359 7572 30393
rect 7740 30359 7756 30393
rect 7556 30321 7756 30359
rect 7814 30393 8014 30409
rect 7814 30359 7830 30393
rect 7998 30359 8014 30393
rect 7814 30321 8014 30359
rect 8072 30393 8272 30409
rect 8072 30359 8088 30393
rect 8256 30359 8272 30393
rect 8072 30321 8272 30359
rect 8330 30393 8530 30409
rect 8330 30359 8346 30393
rect 8514 30359 8530 30393
rect 8330 30321 8530 30359
rect 8588 30393 8788 30409
rect 8588 30359 8604 30393
rect 8772 30359 8788 30393
rect 8588 30321 8788 30359
rect 8846 30393 9046 30409
rect 8846 30359 8862 30393
rect 9030 30359 9046 30393
rect 8846 30321 9046 30359
rect 9104 30393 9304 30409
rect 9104 30359 9120 30393
rect 9288 30359 9304 30393
rect 9104 30321 9304 30359
rect 9362 30393 9562 30409
rect 9362 30359 9378 30393
rect 9546 30359 9562 30393
rect 9362 30321 9562 30359
rect 9620 30393 9820 30409
rect 9620 30359 9636 30393
rect 9804 30359 9820 30393
rect 9620 30321 9820 30359
rect 9878 30393 10078 30409
rect 9878 30359 9894 30393
rect 10062 30359 10078 30393
rect 9878 30321 10078 30359
rect 10136 30393 10336 30409
rect 10136 30359 10152 30393
rect 10320 30359 10336 30393
rect 10136 30321 10336 30359
rect 10394 30393 10594 30409
rect 10394 30359 10410 30393
rect 10578 30359 10594 30393
rect 10394 30321 10594 30359
rect 7556 30211 7756 30237
rect 7814 30211 8014 30237
rect 8072 30211 8272 30237
rect 8330 30211 8530 30237
rect 8588 30211 8788 30237
rect 8846 30211 9046 30237
rect 9104 30211 9304 30237
rect 9362 30211 9562 30237
rect 9620 30211 9820 30237
rect 9878 30211 10078 30237
rect 10136 30211 10336 30237
rect 10394 30211 10594 30237
rect 12939 31889 13139 31915
rect 13197 31889 13397 31915
rect 12939 31651 13139 31689
rect 12939 31617 12955 31651
rect 13123 31617 13139 31651
rect 12939 31601 13139 31617
rect 13197 31651 13397 31689
rect 13197 31617 13213 31651
rect 13381 31617 13397 31651
rect 13197 31601 13397 31617
rect 12939 31006 13139 31022
rect 12939 30972 12955 31006
rect 13123 30972 13139 31006
rect 12939 30925 13139 30972
rect 13197 31006 13397 31022
rect 13197 30972 13213 31006
rect 13381 30972 13397 31006
rect 13197 30925 13397 30972
rect 12939 30699 13139 30725
rect 13197 30699 13397 30725
rect 12939 30429 13139 30455
rect 13197 30429 13397 30455
rect 12939 30191 13139 30229
rect 12939 30157 12955 30191
rect 13123 30157 13139 30191
rect 12939 30141 13139 30157
rect 13197 30191 13397 30229
rect 13197 30157 13213 30191
rect 13381 30157 13397 30191
rect 13197 30141 13397 30157
rect 12686 29477 12716 29503
rect 12770 29477 12800 29503
rect 12854 29477 12884 29503
rect 12938 29477 12968 29503
rect 13022 29477 13052 29503
rect 13106 29477 13136 29503
rect 13190 29477 13220 29503
rect 13274 29477 13304 29503
rect 20288 31108 20488 31134
rect 20546 31108 20746 31134
rect 20804 31108 21004 31134
rect 21062 31108 21262 31134
rect 21320 31108 21520 31134
rect 21578 31108 21778 31134
rect 21836 31108 22036 31134
rect 22094 31108 22294 31134
rect 22352 31108 22552 31134
rect 22610 31108 22810 31134
rect 22868 31108 23068 31134
rect 23126 31108 23326 31134
rect 20288 30861 20488 30908
rect 20288 30827 20304 30861
rect 20472 30827 20488 30861
rect 20288 30811 20488 30827
rect 20546 30861 20746 30908
rect 20546 30827 20562 30861
rect 20730 30827 20746 30861
rect 20546 30811 20746 30827
rect 20804 30861 21004 30908
rect 20804 30827 20820 30861
rect 20988 30827 21004 30861
rect 20804 30811 21004 30827
rect 21062 30861 21262 30908
rect 21062 30827 21078 30861
rect 21246 30827 21262 30861
rect 21062 30811 21262 30827
rect 21320 30861 21520 30908
rect 21320 30827 21336 30861
rect 21504 30827 21520 30861
rect 21320 30811 21520 30827
rect 21578 30861 21778 30908
rect 21578 30827 21594 30861
rect 21762 30827 21778 30861
rect 21578 30811 21778 30827
rect 21836 30861 22036 30908
rect 21836 30827 21852 30861
rect 22020 30827 22036 30861
rect 21836 30811 22036 30827
rect 22094 30861 22294 30908
rect 22094 30827 22110 30861
rect 22278 30827 22294 30861
rect 22094 30811 22294 30827
rect 22352 30861 22552 30908
rect 22352 30827 22368 30861
rect 22536 30827 22552 30861
rect 22352 30811 22552 30827
rect 22610 30861 22810 30908
rect 22610 30827 22626 30861
rect 22794 30827 22810 30861
rect 22610 30811 22810 30827
rect 22868 30861 23068 30908
rect 22868 30827 22884 30861
rect 23052 30827 23068 30861
rect 22868 30811 23068 30827
rect 23126 30861 23326 30908
rect 23126 30827 23142 30861
rect 23310 30827 23326 30861
rect 23126 30811 23326 30827
rect 20546 30753 20746 30769
rect 20546 30719 20562 30753
rect 20730 30719 20746 30753
rect 20288 30681 20488 30707
rect 20546 30681 20746 30719
rect 21320 30753 21520 30769
rect 21320 30719 21336 30753
rect 21504 30719 21520 30753
rect 20804 30681 21004 30707
rect 21062 30681 21262 30707
rect 21320 30681 21520 30719
rect 21578 30753 21778 30769
rect 21578 30719 21594 30753
rect 21762 30719 21778 30753
rect 21578 30681 21778 30719
rect 22352 30753 22552 30769
rect 22352 30719 22368 30753
rect 22536 30719 22552 30753
rect 21836 30681 22036 30707
rect 22094 30681 22294 30707
rect 22352 30681 22552 30719
rect 22610 30753 22810 30769
rect 22610 30719 22626 30753
rect 22794 30719 22810 30753
rect 22610 30681 22810 30719
rect 22868 30681 23068 30707
rect 23126 30681 23326 30707
rect 20288 30443 20488 30481
rect 20546 30455 20746 30481
rect 20288 30409 20304 30443
rect 20472 30409 20488 30443
rect 20288 30393 20488 30409
rect 20804 30443 21004 30481
rect 20804 30409 20820 30443
rect 20988 30409 21004 30443
rect 20804 30393 21004 30409
rect 21062 30443 21262 30481
rect 21320 30455 21520 30481
rect 21578 30455 21778 30481
rect 21062 30409 21078 30443
rect 21246 30409 21262 30443
rect 21062 30393 21262 30409
rect 21836 30443 22036 30481
rect 21836 30409 21852 30443
rect 22020 30409 22036 30443
rect 21836 30393 22036 30409
rect 22094 30443 22294 30481
rect 22352 30455 22552 30481
rect 22610 30455 22810 30481
rect 22094 30409 22110 30443
rect 22278 30409 22294 30443
rect 22094 30393 22294 30409
rect 22868 30443 23068 30481
rect 22868 30409 22884 30443
rect 23052 30409 23068 30443
rect 22868 30393 23068 30409
rect 23126 30443 23326 30481
rect 23126 30409 23142 30443
rect 23310 30409 23326 30443
rect 23126 30393 23326 30409
rect 20288 30317 20488 30333
rect 20288 30283 20304 30317
rect 20472 30283 20488 30317
rect 20288 30245 20488 30283
rect 20546 30317 20746 30333
rect 20546 30283 20562 30317
rect 20730 30283 20746 30317
rect 20546 30245 20746 30283
rect 20804 30317 21004 30333
rect 20804 30283 20820 30317
rect 20988 30283 21004 30317
rect 20804 30245 21004 30283
rect 21062 30317 21262 30333
rect 21062 30283 21078 30317
rect 21246 30283 21262 30317
rect 21062 30245 21262 30283
rect 21320 30317 21520 30333
rect 21320 30283 21336 30317
rect 21504 30283 21520 30317
rect 21320 30245 21520 30283
rect 21578 30317 21778 30333
rect 21578 30283 21594 30317
rect 21762 30283 21778 30317
rect 21578 30245 21778 30283
rect 21836 30317 22036 30333
rect 21836 30283 21852 30317
rect 22020 30283 22036 30317
rect 21836 30245 22036 30283
rect 22094 30317 22294 30333
rect 22094 30283 22110 30317
rect 22278 30283 22294 30317
rect 22094 30245 22294 30283
rect 22352 30317 22552 30333
rect 22352 30283 22368 30317
rect 22536 30283 22552 30317
rect 22352 30245 22552 30283
rect 22610 30317 22810 30333
rect 22610 30283 22626 30317
rect 22794 30283 22810 30317
rect 22610 30245 22810 30283
rect 22868 30317 23068 30333
rect 22868 30283 22884 30317
rect 23052 30283 23068 30317
rect 22868 30245 23068 30283
rect 23126 30317 23326 30333
rect 23126 30283 23142 30317
rect 23310 30283 23326 30317
rect 23126 30245 23326 30283
rect 20288 30135 20488 30161
rect 20546 30135 20746 30161
rect 20804 30135 21004 30161
rect 21062 30135 21262 30161
rect 21320 30135 21520 30161
rect 21578 30135 21778 30161
rect 21836 30135 22036 30161
rect 22094 30135 22294 30161
rect 22352 30135 22552 30161
rect 22610 30135 22810 30161
rect 22868 30135 23068 30161
rect 23126 30135 23326 30161
rect 12686 29245 12716 29277
rect 12770 29245 12800 29277
rect 12854 29245 12884 29277
rect 12938 29245 12968 29277
rect 13022 29245 13052 29277
rect 13106 29245 13136 29277
rect 13190 29245 13220 29277
rect 13274 29245 13304 29277
rect 12686 29229 13304 29245
rect 12686 29195 12726 29229
rect 12760 29195 12810 29229
rect 12844 29195 12894 29229
rect 12928 29195 12978 29229
rect 13012 29195 13062 29229
rect 13096 29195 13146 29229
rect 13180 29195 13230 29229
rect 13264 29195 13304 29229
rect 12686 29179 13304 29195
rect 12686 29157 12716 29179
rect 12770 29157 12800 29179
rect 12854 29157 12884 29179
rect 12938 29157 12968 29179
rect 13022 29157 13052 29179
rect 13106 29157 13136 29179
rect 13190 29157 13220 29179
rect 13274 29157 13304 29179
rect 12686 29001 12716 29027
rect 12770 29001 12800 29027
rect 12854 29001 12884 29027
rect 12938 29001 12968 29027
rect 13022 29001 13052 29027
rect 13106 29001 13136 29027
rect 13190 29001 13220 29027
rect 13274 29001 13304 29027
rect 25671 31813 25871 31839
rect 25929 31813 26129 31839
rect 25671 31575 25871 31613
rect 25671 31541 25687 31575
rect 25855 31541 25871 31575
rect 25671 31525 25871 31541
rect 25929 31575 26129 31613
rect 25929 31541 25945 31575
rect 26113 31541 26129 31575
rect 25929 31525 26129 31541
rect 25671 30930 25871 30946
rect 25671 30896 25687 30930
rect 25855 30896 25871 30930
rect 25671 30849 25871 30896
rect 25929 30930 26129 30946
rect 25929 30896 25945 30930
rect 26113 30896 26129 30930
rect 25929 30849 26129 30896
rect 25671 30623 25871 30649
rect 25929 30623 26129 30649
rect 25671 30353 25871 30379
rect 25929 30353 26129 30379
rect 25671 30115 25871 30153
rect 25671 30081 25687 30115
rect 25855 30081 25871 30115
rect 25671 30065 25871 30081
rect 25929 30115 26129 30153
rect 25929 30081 25945 30115
rect 26113 30081 26129 30115
rect 25929 30065 26129 30081
rect 25418 29401 25448 29427
rect 25502 29401 25532 29427
rect 25586 29401 25616 29427
rect 25670 29401 25700 29427
rect 25754 29401 25784 29427
rect 25838 29401 25868 29427
rect 25922 29401 25952 29427
rect 26006 29401 26036 29427
rect 25418 29169 25448 29201
rect 25502 29169 25532 29201
rect 25586 29169 25616 29201
rect 25670 29169 25700 29201
rect 25754 29169 25784 29201
rect 25838 29169 25868 29201
rect 25922 29169 25952 29201
rect 26006 29169 26036 29201
rect 25418 29153 26036 29169
rect 25418 29119 25458 29153
rect 25492 29119 25542 29153
rect 25576 29119 25626 29153
rect 25660 29119 25710 29153
rect 25744 29119 25794 29153
rect 25828 29119 25878 29153
rect 25912 29119 25962 29153
rect 25996 29119 26036 29153
rect 25418 29103 26036 29119
rect 25418 29081 25448 29103
rect 25502 29081 25532 29103
rect 25586 29081 25616 29103
rect 25670 29081 25700 29103
rect 25754 29081 25784 29103
rect 25838 29081 25868 29103
rect 25922 29081 25952 29103
rect 26006 29081 26036 29103
rect 25418 28925 25448 28951
rect 25502 28925 25532 28951
rect 25586 28925 25616 28951
rect 25670 28925 25700 28951
rect 25754 28925 25784 28951
rect 25838 28925 25868 28951
rect 25922 28925 25952 28951
rect 26006 28925 26036 28951
rect 13059 25762 13259 25778
rect 13059 25728 13075 25762
rect 13243 25728 13259 25762
rect 13059 25681 13259 25728
rect 13317 25762 13517 25778
rect 13317 25728 13333 25762
rect 13501 25728 13517 25762
rect 13317 25681 13517 25728
rect 13059 25455 13259 25481
rect 13317 25455 13517 25481
rect 25767 25632 25967 25648
rect 25767 25598 25783 25632
rect 25951 25598 25967 25632
rect 25767 25551 25967 25598
rect 26025 25632 26225 25648
rect 26025 25598 26041 25632
rect 26209 25598 26225 25632
rect 26025 25551 26225 25598
rect 7676 24480 7876 24506
rect 7934 24480 8134 24506
rect 8192 24480 8392 24506
rect 8450 24480 8650 24506
rect 8708 24480 8908 24506
rect 8966 24480 9166 24506
rect 9224 24480 9424 24506
rect 9482 24480 9682 24506
rect 9740 24480 9940 24506
rect 9998 24480 10198 24506
rect 10256 24480 10456 24506
rect 10514 24480 10714 24506
rect 7676 24233 7876 24280
rect 7676 24199 7692 24233
rect 7860 24199 7876 24233
rect 7676 24183 7876 24199
rect 7934 24233 8134 24280
rect 7934 24199 7950 24233
rect 8118 24199 8134 24233
rect 7934 24183 8134 24199
rect 8192 24233 8392 24280
rect 8192 24199 8208 24233
rect 8376 24199 8392 24233
rect 8192 24183 8392 24199
rect 8450 24233 8650 24280
rect 8450 24199 8466 24233
rect 8634 24199 8650 24233
rect 8450 24183 8650 24199
rect 8708 24233 8908 24280
rect 8708 24199 8724 24233
rect 8892 24199 8908 24233
rect 8708 24183 8908 24199
rect 8966 24233 9166 24280
rect 8966 24199 8982 24233
rect 9150 24199 9166 24233
rect 8966 24183 9166 24199
rect 9224 24233 9424 24280
rect 9224 24199 9240 24233
rect 9408 24199 9424 24233
rect 9224 24183 9424 24199
rect 9482 24233 9682 24280
rect 9482 24199 9498 24233
rect 9666 24199 9682 24233
rect 9482 24183 9682 24199
rect 9740 24233 9940 24280
rect 9740 24199 9756 24233
rect 9924 24199 9940 24233
rect 9740 24183 9940 24199
rect 9998 24233 10198 24280
rect 9998 24199 10014 24233
rect 10182 24199 10198 24233
rect 9998 24183 10198 24199
rect 10256 24233 10456 24280
rect 10256 24199 10272 24233
rect 10440 24199 10456 24233
rect 10256 24183 10456 24199
rect 10514 24233 10714 24280
rect 10514 24199 10530 24233
rect 10698 24199 10714 24233
rect 10514 24183 10714 24199
rect 7934 24125 8134 24141
rect 7934 24091 7950 24125
rect 8118 24091 8134 24125
rect 7676 24053 7876 24079
rect 7934 24053 8134 24091
rect 8708 24125 8908 24141
rect 8708 24091 8724 24125
rect 8892 24091 8908 24125
rect 8192 24053 8392 24079
rect 8450 24053 8650 24079
rect 8708 24053 8908 24091
rect 8966 24125 9166 24141
rect 8966 24091 8982 24125
rect 9150 24091 9166 24125
rect 8966 24053 9166 24091
rect 9740 24125 9940 24141
rect 9740 24091 9756 24125
rect 9924 24091 9940 24125
rect 9224 24053 9424 24079
rect 9482 24053 9682 24079
rect 9740 24053 9940 24091
rect 9998 24125 10198 24141
rect 9998 24091 10014 24125
rect 10182 24091 10198 24125
rect 9998 24053 10198 24091
rect 10256 24053 10456 24079
rect 10514 24053 10714 24079
rect 7676 23815 7876 23853
rect 7934 23827 8134 23853
rect 7676 23781 7692 23815
rect 7860 23781 7876 23815
rect 7676 23765 7876 23781
rect 8192 23815 8392 23853
rect 8192 23781 8208 23815
rect 8376 23781 8392 23815
rect 8192 23765 8392 23781
rect 8450 23815 8650 23853
rect 8708 23827 8908 23853
rect 8966 23827 9166 23853
rect 8450 23781 8466 23815
rect 8634 23781 8650 23815
rect 8450 23765 8650 23781
rect 9224 23815 9424 23853
rect 9224 23781 9240 23815
rect 9408 23781 9424 23815
rect 9224 23765 9424 23781
rect 9482 23815 9682 23853
rect 9740 23827 9940 23853
rect 9998 23827 10198 23853
rect 9482 23781 9498 23815
rect 9666 23781 9682 23815
rect 9482 23765 9682 23781
rect 10256 23815 10456 23853
rect 10256 23781 10272 23815
rect 10440 23781 10456 23815
rect 10256 23765 10456 23781
rect 10514 23815 10714 23853
rect 10514 23781 10530 23815
rect 10698 23781 10714 23815
rect 10514 23765 10714 23781
rect 7676 23689 7876 23705
rect 7676 23655 7692 23689
rect 7860 23655 7876 23689
rect 7676 23617 7876 23655
rect 7934 23689 8134 23705
rect 7934 23655 7950 23689
rect 8118 23655 8134 23689
rect 7934 23617 8134 23655
rect 8192 23689 8392 23705
rect 8192 23655 8208 23689
rect 8376 23655 8392 23689
rect 8192 23617 8392 23655
rect 8450 23689 8650 23705
rect 8450 23655 8466 23689
rect 8634 23655 8650 23689
rect 8450 23617 8650 23655
rect 8708 23689 8908 23705
rect 8708 23655 8724 23689
rect 8892 23655 8908 23689
rect 8708 23617 8908 23655
rect 8966 23689 9166 23705
rect 8966 23655 8982 23689
rect 9150 23655 9166 23689
rect 8966 23617 9166 23655
rect 9224 23689 9424 23705
rect 9224 23655 9240 23689
rect 9408 23655 9424 23689
rect 9224 23617 9424 23655
rect 9482 23689 9682 23705
rect 9482 23655 9498 23689
rect 9666 23655 9682 23689
rect 9482 23617 9682 23655
rect 9740 23689 9940 23705
rect 9740 23655 9756 23689
rect 9924 23655 9940 23689
rect 9740 23617 9940 23655
rect 9998 23689 10198 23705
rect 9998 23655 10014 23689
rect 10182 23655 10198 23689
rect 9998 23617 10198 23655
rect 10256 23689 10456 23705
rect 10256 23655 10272 23689
rect 10440 23655 10456 23689
rect 10256 23617 10456 23655
rect 10514 23689 10714 23705
rect 10514 23655 10530 23689
rect 10698 23655 10714 23689
rect 10514 23617 10714 23655
rect 7676 23507 7876 23533
rect 7934 23507 8134 23533
rect 8192 23507 8392 23533
rect 8450 23507 8650 23533
rect 8708 23507 8908 23533
rect 8966 23507 9166 23533
rect 9224 23507 9424 23533
rect 9482 23507 9682 23533
rect 9740 23507 9940 23533
rect 9998 23507 10198 23533
rect 10256 23507 10456 23533
rect 10514 23507 10714 23533
rect 13059 25185 13259 25211
rect 13317 25185 13517 25211
rect 25767 25325 25967 25351
rect 26025 25325 26225 25351
rect 13059 24947 13259 24985
rect 13059 24913 13075 24947
rect 13243 24913 13259 24947
rect 13059 24897 13259 24913
rect 13317 24947 13517 24985
rect 13317 24913 13333 24947
rect 13501 24913 13517 24947
rect 13317 24897 13517 24913
rect 13059 24302 13259 24318
rect 13059 24268 13075 24302
rect 13243 24268 13259 24302
rect 13059 24221 13259 24268
rect 13317 24302 13517 24318
rect 13317 24268 13333 24302
rect 13501 24268 13517 24302
rect 13317 24221 13517 24268
rect 13059 23995 13259 24021
rect 13317 23995 13517 24021
rect 13059 23725 13259 23751
rect 13317 23725 13517 23751
rect 13059 23487 13259 23525
rect 13059 23453 13075 23487
rect 13243 23453 13259 23487
rect 13059 23437 13259 23453
rect 13317 23487 13517 23525
rect 13317 23453 13333 23487
rect 13501 23453 13517 23487
rect 13317 23437 13517 23453
rect 12806 22773 12836 22799
rect 12890 22773 12920 22799
rect 12974 22773 13004 22799
rect 13058 22773 13088 22799
rect 13142 22773 13172 22799
rect 13226 22773 13256 22799
rect 13310 22773 13340 22799
rect 13394 22773 13424 22799
rect 12806 22541 12836 22573
rect 12890 22541 12920 22573
rect 12974 22541 13004 22573
rect 13058 22541 13088 22573
rect 13142 22541 13172 22573
rect 13226 22541 13256 22573
rect 13310 22541 13340 22573
rect 13394 22541 13424 22573
rect 12806 22525 13424 22541
rect 12806 22491 12846 22525
rect 12880 22491 12930 22525
rect 12964 22491 13014 22525
rect 13048 22491 13098 22525
rect 13132 22491 13182 22525
rect 13216 22491 13266 22525
rect 13300 22491 13350 22525
rect 13384 22491 13424 22525
rect 12806 22475 13424 22491
rect 20384 24350 20584 24376
rect 20642 24350 20842 24376
rect 20900 24350 21100 24376
rect 21158 24350 21358 24376
rect 21416 24350 21616 24376
rect 21674 24350 21874 24376
rect 21932 24350 22132 24376
rect 22190 24350 22390 24376
rect 22448 24350 22648 24376
rect 22706 24350 22906 24376
rect 22964 24350 23164 24376
rect 23222 24350 23422 24376
rect 20384 24103 20584 24150
rect 20384 24069 20400 24103
rect 20568 24069 20584 24103
rect 20384 24053 20584 24069
rect 20642 24103 20842 24150
rect 20642 24069 20658 24103
rect 20826 24069 20842 24103
rect 20642 24053 20842 24069
rect 20900 24103 21100 24150
rect 20900 24069 20916 24103
rect 21084 24069 21100 24103
rect 20900 24053 21100 24069
rect 21158 24103 21358 24150
rect 21158 24069 21174 24103
rect 21342 24069 21358 24103
rect 21158 24053 21358 24069
rect 21416 24103 21616 24150
rect 21416 24069 21432 24103
rect 21600 24069 21616 24103
rect 21416 24053 21616 24069
rect 21674 24103 21874 24150
rect 21674 24069 21690 24103
rect 21858 24069 21874 24103
rect 21674 24053 21874 24069
rect 21932 24103 22132 24150
rect 21932 24069 21948 24103
rect 22116 24069 22132 24103
rect 21932 24053 22132 24069
rect 22190 24103 22390 24150
rect 22190 24069 22206 24103
rect 22374 24069 22390 24103
rect 22190 24053 22390 24069
rect 22448 24103 22648 24150
rect 22448 24069 22464 24103
rect 22632 24069 22648 24103
rect 22448 24053 22648 24069
rect 22706 24103 22906 24150
rect 22706 24069 22722 24103
rect 22890 24069 22906 24103
rect 22706 24053 22906 24069
rect 22964 24103 23164 24150
rect 22964 24069 22980 24103
rect 23148 24069 23164 24103
rect 22964 24053 23164 24069
rect 23222 24103 23422 24150
rect 23222 24069 23238 24103
rect 23406 24069 23422 24103
rect 23222 24053 23422 24069
rect 20642 23995 20842 24011
rect 20642 23961 20658 23995
rect 20826 23961 20842 23995
rect 20384 23923 20584 23949
rect 20642 23923 20842 23961
rect 21416 23995 21616 24011
rect 21416 23961 21432 23995
rect 21600 23961 21616 23995
rect 20900 23923 21100 23949
rect 21158 23923 21358 23949
rect 21416 23923 21616 23961
rect 21674 23995 21874 24011
rect 21674 23961 21690 23995
rect 21858 23961 21874 23995
rect 21674 23923 21874 23961
rect 22448 23995 22648 24011
rect 22448 23961 22464 23995
rect 22632 23961 22648 23995
rect 21932 23923 22132 23949
rect 22190 23923 22390 23949
rect 22448 23923 22648 23961
rect 22706 23995 22906 24011
rect 22706 23961 22722 23995
rect 22890 23961 22906 23995
rect 22706 23923 22906 23961
rect 22964 23923 23164 23949
rect 23222 23923 23422 23949
rect 20384 23685 20584 23723
rect 20642 23697 20842 23723
rect 20384 23651 20400 23685
rect 20568 23651 20584 23685
rect 20384 23635 20584 23651
rect 20900 23685 21100 23723
rect 20900 23651 20916 23685
rect 21084 23651 21100 23685
rect 20900 23635 21100 23651
rect 21158 23685 21358 23723
rect 21416 23697 21616 23723
rect 21674 23697 21874 23723
rect 21158 23651 21174 23685
rect 21342 23651 21358 23685
rect 21158 23635 21358 23651
rect 21932 23685 22132 23723
rect 21932 23651 21948 23685
rect 22116 23651 22132 23685
rect 21932 23635 22132 23651
rect 22190 23685 22390 23723
rect 22448 23697 22648 23723
rect 22706 23697 22906 23723
rect 22190 23651 22206 23685
rect 22374 23651 22390 23685
rect 22190 23635 22390 23651
rect 22964 23685 23164 23723
rect 22964 23651 22980 23685
rect 23148 23651 23164 23685
rect 22964 23635 23164 23651
rect 23222 23685 23422 23723
rect 23222 23651 23238 23685
rect 23406 23651 23422 23685
rect 23222 23635 23422 23651
rect 20384 23559 20584 23575
rect 20384 23525 20400 23559
rect 20568 23525 20584 23559
rect 20384 23487 20584 23525
rect 20642 23559 20842 23575
rect 20642 23525 20658 23559
rect 20826 23525 20842 23559
rect 20642 23487 20842 23525
rect 20900 23559 21100 23575
rect 20900 23525 20916 23559
rect 21084 23525 21100 23559
rect 20900 23487 21100 23525
rect 21158 23559 21358 23575
rect 21158 23525 21174 23559
rect 21342 23525 21358 23559
rect 21158 23487 21358 23525
rect 21416 23559 21616 23575
rect 21416 23525 21432 23559
rect 21600 23525 21616 23559
rect 21416 23487 21616 23525
rect 21674 23559 21874 23575
rect 21674 23525 21690 23559
rect 21858 23525 21874 23559
rect 21674 23487 21874 23525
rect 21932 23559 22132 23575
rect 21932 23525 21948 23559
rect 22116 23525 22132 23559
rect 21932 23487 22132 23525
rect 22190 23559 22390 23575
rect 22190 23525 22206 23559
rect 22374 23525 22390 23559
rect 22190 23487 22390 23525
rect 22448 23559 22648 23575
rect 22448 23525 22464 23559
rect 22632 23525 22648 23559
rect 22448 23487 22648 23525
rect 22706 23559 22906 23575
rect 22706 23525 22722 23559
rect 22890 23525 22906 23559
rect 22706 23487 22906 23525
rect 22964 23559 23164 23575
rect 22964 23525 22980 23559
rect 23148 23525 23164 23559
rect 22964 23487 23164 23525
rect 23222 23559 23422 23575
rect 23222 23525 23238 23559
rect 23406 23525 23422 23559
rect 23222 23487 23422 23525
rect 20384 23377 20584 23403
rect 20642 23377 20842 23403
rect 20900 23377 21100 23403
rect 21158 23377 21358 23403
rect 21416 23377 21616 23403
rect 21674 23377 21874 23403
rect 21932 23377 22132 23403
rect 22190 23377 22390 23403
rect 22448 23377 22648 23403
rect 22706 23377 22906 23403
rect 22964 23377 23164 23403
rect 23222 23377 23422 23403
rect 12806 22453 12836 22475
rect 12890 22453 12920 22475
rect 12974 22453 13004 22475
rect 13058 22453 13088 22475
rect 13142 22453 13172 22475
rect 13226 22453 13256 22475
rect 13310 22453 13340 22475
rect 13394 22453 13424 22475
rect 12806 22297 12836 22323
rect 12890 22297 12920 22323
rect 12974 22297 13004 22323
rect 13058 22297 13088 22323
rect 13142 22297 13172 22323
rect 13226 22297 13256 22323
rect 13310 22297 13340 22323
rect 13394 22297 13424 22323
rect 25767 25055 25967 25081
rect 26025 25055 26225 25081
rect 25767 24817 25967 24855
rect 25767 24783 25783 24817
rect 25951 24783 25967 24817
rect 25767 24767 25967 24783
rect 26025 24817 26225 24855
rect 26025 24783 26041 24817
rect 26209 24783 26225 24817
rect 26025 24767 26225 24783
rect 25767 24172 25967 24188
rect 25767 24138 25783 24172
rect 25951 24138 25967 24172
rect 25767 24091 25967 24138
rect 26025 24172 26225 24188
rect 26025 24138 26041 24172
rect 26209 24138 26225 24172
rect 26025 24091 26225 24138
rect 25767 23865 25967 23891
rect 26025 23865 26225 23891
rect 25767 23595 25967 23621
rect 26025 23595 26225 23621
rect 25767 23357 25967 23395
rect 25767 23323 25783 23357
rect 25951 23323 25967 23357
rect 25767 23307 25967 23323
rect 26025 23357 26225 23395
rect 26025 23323 26041 23357
rect 26209 23323 26225 23357
rect 26025 23307 26225 23323
rect 25514 22643 25544 22669
rect 25598 22643 25628 22669
rect 25682 22643 25712 22669
rect 25766 22643 25796 22669
rect 25850 22643 25880 22669
rect 25934 22643 25964 22669
rect 26018 22643 26048 22669
rect 26102 22643 26132 22669
rect 25514 22411 25544 22443
rect 25598 22411 25628 22443
rect 25682 22411 25712 22443
rect 25766 22411 25796 22443
rect 25850 22411 25880 22443
rect 25934 22411 25964 22443
rect 26018 22411 26048 22443
rect 26102 22411 26132 22443
rect 25514 22395 26132 22411
rect 25514 22361 25554 22395
rect 25588 22361 25638 22395
rect 25672 22361 25722 22395
rect 25756 22361 25806 22395
rect 25840 22361 25890 22395
rect 25924 22361 25974 22395
rect 26008 22361 26058 22395
rect 26092 22361 26132 22395
rect 25514 22345 26132 22361
rect 25514 22323 25544 22345
rect 25598 22323 25628 22345
rect 25682 22323 25712 22345
rect 25766 22323 25796 22345
rect 25850 22323 25880 22345
rect 25934 22323 25964 22345
rect 26018 22323 26048 22345
rect 26102 22323 26132 22345
rect 25514 22167 25544 22193
rect 25598 22167 25628 22193
rect 25682 22167 25712 22193
rect 25766 22167 25796 22193
rect 25850 22167 25880 22193
rect 25934 22167 25964 22193
rect 26018 22167 26048 22193
rect 26102 22167 26132 22193
rect 12935 18716 13135 18732
rect 12935 18682 12951 18716
rect 13119 18682 13135 18716
rect 12935 18635 13135 18682
rect 13193 18716 13393 18732
rect 13193 18682 13209 18716
rect 13377 18682 13393 18716
rect 13193 18635 13393 18682
rect 12935 18409 13135 18435
rect 13193 18409 13393 18435
rect 26117 18586 26317 18602
rect 26117 18552 26133 18586
rect 26301 18552 26317 18586
rect 26117 18505 26317 18552
rect 26375 18586 26575 18602
rect 26375 18552 26391 18586
rect 26559 18552 26575 18586
rect 26375 18505 26575 18552
rect 7552 17434 7752 17460
rect 7810 17434 8010 17460
rect 8068 17434 8268 17460
rect 8326 17434 8526 17460
rect 8584 17434 8784 17460
rect 8842 17434 9042 17460
rect 9100 17434 9300 17460
rect 9358 17434 9558 17460
rect 9616 17434 9816 17460
rect 9874 17434 10074 17460
rect 10132 17434 10332 17460
rect 10390 17434 10590 17460
rect 7552 17187 7752 17234
rect 7552 17153 7568 17187
rect 7736 17153 7752 17187
rect 7552 17137 7752 17153
rect 7810 17187 8010 17234
rect 7810 17153 7826 17187
rect 7994 17153 8010 17187
rect 7810 17137 8010 17153
rect 8068 17187 8268 17234
rect 8068 17153 8084 17187
rect 8252 17153 8268 17187
rect 8068 17137 8268 17153
rect 8326 17187 8526 17234
rect 8326 17153 8342 17187
rect 8510 17153 8526 17187
rect 8326 17137 8526 17153
rect 8584 17187 8784 17234
rect 8584 17153 8600 17187
rect 8768 17153 8784 17187
rect 8584 17137 8784 17153
rect 8842 17187 9042 17234
rect 8842 17153 8858 17187
rect 9026 17153 9042 17187
rect 8842 17137 9042 17153
rect 9100 17187 9300 17234
rect 9100 17153 9116 17187
rect 9284 17153 9300 17187
rect 9100 17137 9300 17153
rect 9358 17187 9558 17234
rect 9358 17153 9374 17187
rect 9542 17153 9558 17187
rect 9358 17137 9558 17153
rect 9616 17187 9816 17234
rect 9616 17153 9632 17187
rect 9800 17153 9816 17187
rect 9616 17137 9816 17153
rect 9874 17187 10074 17234
rect 9874 17153 9890 17187
rect 10058 17153 10074 17187
rect 9874 17137 10074 17153
rect 10132 17187 10332 17234
rect 10132 17153 10148 17187
rect 10316 17153 10332 17187
rect 10132 17137 10332 17153
rect 10390 17187 10590 17234
rect 10390 17153 10406 17187
rect 10574 17153 10590 17187
rect 10390 17137 10590 17153
rect 7810 17079 8010 17095
rect 7810 17045 7826 17079
rect 7994 17045 8010 17079
rect 7552 17007 7752 17033
rect 7810 17007 8010 17045
rect 8584 17079 8784 17095
rect 8584 17045 8600 17079
rect 8768 17045 8784 17079
rect 8068 17007 8268 17033
rect 8326 17007 8526 17033
rect 8584 17007 8784 17045
rect 8842 17079 9042 17095
rect 8842 17045 8858 17079
rect 9026 17045 9042 17079
rect 8842 17007 9042 17045
rect 9616 17079 9816 17095
rect 9616 17045 9632 17079
rect 9800 17045 9816 17079
rect 9100 17007 9300 17033
rect 9358 17007 9558 17033
rect 9616 17007 9816 17045
rect 9874 17079 10074 17095
rect 9874 17045 9890 17079
rect 10058 17045 10074 17079
rect 9874 17007 10074 17045
rect 10132 17007 10332 17033
rect 10390 17007 10590 17033
rect 7552 16769 7752 16807
rect 7810 16781 8010 16807
rect 7552 16735 7568 16769
rect 7736 16735 7752 16769
rect 7552 16719 7752 16735
rect 8068 16769 8268 16807
rect 8068 16735 8084 16769
rect 8252 16735 8268 16769
rect 8068 16719 8268 16735
rect 8326 16769 8526 16807
rect 8584 16781 8784 16807
rect 8842 16781 9042 16807
rect 8326 16735 8342 16769
rect 8510 16735 8526 16769
rect 8326 16719 8526 16735
rect 9100 16769 9300 16807
rect 9100 16735 9116 16769
rect 9284 16735 9300 16769
rect 9100 16719 9300 16735
rect 9358 16769 9558 16807
rect 9616 16781 9816 16807
rect 9874 16781 10074 16807
rect 9358 16735 9374 16769
rect 9542 16735 9558 16769
rect 9358 16719 9558 16735
rect 10132 16769 10332 16807
rect 10132 16735 10148 16769
rect 10316 16735 10332 16769
rect 10132 16719 10332 16735
rect 10390 16769 10590 16807
rect 10390 16735 10406 16769
rect 10574 16735 10590 16769
rect 10390 16719 10590 16735
rect 7552 16643 7752 16659
rect 7552 16609 7568 16643
rect 7736 16609 7752 16643
rect 7552 16571 7752 16609
rect 7810 16643 8010 16659
rect 7810 16609 7826 16643
rect 7994 16609 8010 16643
rect 7810 16571 8010 16609
rect 8068 16643 8268 16659
rect 8068 16609 8084 16643
rect 8252 16609 8268 16643
rect 8068 16571 8268 16609
rect 8326 16643 8526 16659
rect 8326 16609 8342 16643
rect 8510 16609 8526 16643
rect 8326 16571 8526 16609
rect 8584 16643 8784 16659
rect 8584 16609 8600 16643
rect 8768 16609 8784 16643
rect 8584 16571 8784 16609
rect 8842 16643 9042 16659
rect 8842 16609 8858 16643
rect 9026 16609 9042 16643
rect 8842 16571 9042 16609
rect 9100 16643 9300 16659
rect 9100 16609 9116 16643
rect 9284 16609 9300 16643
rect 9100 16571 9300 16609
rect 9358 16643 9558 16659
rect 9358 16609 9374 16643
rect 9542 16609 9558 16643
rect 9358 16571 9558 16609
rect 9616 16643 9816 16659
rect 9616 16609 9632 16643
rect 9800 16609 9816 16643
rect 9616 16571 9816 16609
rect 9874 16643 10074 16659
rect 9874 16609 9890 16643
rect 10058 16609 10074 16643
rect 9874 16571 10074 16609
rect 10132 16643 10332 16659
rect 10132 16609 10148 16643
rect 10316 16609 10332 16643
rect 10132 16571 10332 16609
rect 10390 16643 10590 16659
rect 10390 16609 10406 16643
rect 10574 16609 10590 16643
rect 10390 16571 10590 16609
rect 7552 16461 7752 16487
rect 7810 16461 8010 16487
rect 8068 16461 8268 16487
rect 8326 16461 8526 16487
rect 8584 16461 8784 16487
rect 8842 16461 9042 16487
rect 9100 16461 9300 16487
rect 9358 16461 9558 16487
rect 9616 16461 9816 16487
rect 9874 16461 10074 16487
rect 10132 16461 10332 16487
rect 10390 16461 10590 16487
rect 12935 18139 13135 18165
rect 13193 18139 13393 18165
rect 26117 18279 26317 18305
rect 26375 18279 26575 18305
rect 12935 17901 13135 17939
rect 12935 17867 12951 17901
rect 13119 17867 13135 17901
rect 12935 17851 13135 17867
rect 13193 17901 13393 17939
rect 13193 17867 13209 17901
rect 13377 17867 13393 17901
rect 13193 17851 13393 17867
rect 12935 17256 13135 17272
rect 12935 17222 12951 17256
rect 13119 17222 13135 17256
rect 12935 17175 13135 17222
rect 13193 17256 13393 17272
rect 13193 17222 13209 17256
rect 13377 17222 13393 17256
rect 13193 17175 13393 17222
rect 12935 16949 13135 16975
rect 13193 16949 13393 16975
rect 12935 16679 13135 16705
rect 13193 16679 13393 16705
rect 12935 16441 13135 16479
rect 12935 16407 12951 16441
rect 13119 16407 13135 16441
rect 12935 16391 13135 16407
rect 13193 16441 13393 16479
rect 13193 16407 13209 16441
rect 13377 16407 13393 16441
rect 13193 16391 13393 16407
rect 12682 15727 12712 15753
rect 12766 15727 12796 15753
rect 12850 15727 12880 15753
rect 12934 15727 12964 15753
rect 13018 15727 13048 15753
rect 13102 15727 13132 15753
rect 13186 15727 13216 15753
rect 13270 15727 13300 15753
rect 12682 15495 12712 15527
rect 12766 15495 12796 15527
rect 12850 15495 12880 15527
rect 12934 15495 12964 15527
rect 13018 15495 13048 15527
rect 13102 15495 13132 15527
rect 13186 15495 13216 15527
rect 13270 15495 13300 15527
rect 12682 15479 13300 15495
rect 12682 15445 12722 15479
rect 12756 15445 12806 15479
rect 12840 15445 12890 15479
rect 12924 15445 12974 15479
rect 13008 15445 13058 15479
rect 13092 15445 13142 15479
rect 13176 15445 13226 15479
rect 13260 15445 13300 15479
rect 12682 15429 13300 15445
rect 20734 17304 20934 17330
rect 20992 17304 21192 17330
rect 21250 17304 21450 17330
rect 21508 17304 21708 17330
rect 21766 17304 21966 17330
rect 22024 17304 22224 17330
rect 22282 17304 22482 17330
rect 22540 17304 22740 17330
rect 22798 17304 22998 17330
rect 23056 17304 23256 17330
rect 23314 17304 23514 17330
rect 23572 17304 23772 17330
rect 20734 17057 20934 17104
rect 20734 17023 20750 17057
rect 20918 17023 20934 17057
rect 20734 17007 20934 17023
rect 20992 17057 21192 17104
rect 20992 17023 21008 17057
rect 21176 17023 21192 17057
rect 20992 17007 21192 17023
rect 21250 17057 21450 17104
rect 21250 17023 21266 17057
rect 21434 17023 21450 17057
rect 21250 17007 21450 17023
rect 21508 17057 21708 17104
rect 21508 17023 21524 17057
rect 21692 17023 21708 17057
rect 21508 17007 21708 17023
rect 21766 17057 21966 17104
rect 21766 17023 21782 17057
rect 21950 17023 21966 17057
rect 21766 17007 21966 17023
rect 22024 17057 22224 17104
rect 22024 17023 22040 17057
rect 22208 17023 22224 17057
rect 22024 17007 22224 17023
rect 22282 17057 22482 17104
rect 22282 17023 22298 17057
rect 22466 17023 22482 17057
rect 22282 17007 22482 17023
rect 22540 17057 22740 17104
rect 22540 17023 22556 17057
rect 22724 17023 22740 17057
rect 22540 17007 22740 17023
rect 22798 17057 22998 17104
rect 22798 17023 22814 17057
rect 22982 17023 22998 17057
rect 22798 17007 22998 17023
rect 23056 17057 23256 17104
rect 23056 17023 23072 17057
rect 23240 17023 23256 17057
rect 23056 17007 23256 17023
rect 23314 17057 23514 17104
rect 23314 17023 23330 17057
rect 23498 17023 23514 17057
rect 23314 17007 23514 17023
rect 23572 17057 23772 17104
rect 23572 17023 23588 17057
rect 23756 17023 23772 17057
rect 23572 17007 23772 17023
rect 20992 16949 21192 16965
rect 20992 16915 21008 16949
rect 21176 16915 21192 16949
rect 20734 16877 20934 16903
rect 20992 16877 21192 16915
rect 21766 16949 21966 16965
rect 21766 16915 21782 16949
rect 21950 16915 21966 16949
rect 21250 16877 21450 16903
rect 21508 16877 21708 16903
rect 21766 16877 21966 16915
rect 22024 16949 22224 16965
rect 22024 16915 22040 16949
rect 22208 16915 22224 16949
rect 22024 16877 22224 16915
rect 22798 16949 22998 16965
rect 22798 16915 22814 16949
rect 22982 16915 22998 16949
rect 22282 16877 22482 16903
rect 22540 16877 22740 16903
rect 22798 16877 22998 16915
rect 23056 16949 23256 16965
rect 23056 16915 23072 16949
rect 23240 16915 23256 16949
rect 23056 16877 23256 16915
rect 23314 16877 23514 16903
rect 23572 16877 23772 16903
rect 20734 16639 20934 16677
rect 20992 16651 21192 16677
rect 20734 16605 20750 16639
rect 20918 16605 20934 16639
rect 20734 16589 20934 16605
rect 21250 16639 21450 16677
rect 21250 16605 21266 16639
rect 21434 16605 21450 16639
rect 21250 16589 21450 16605
rect 21508 16639 21708 16677
rect 21766 16651 21966 16677
rect 22024 16651 22224 16677
rect 21508 16605 21524 16639
rect 21692 16605 21708 16639
rect 21508 16589 21708 16605
rect 22282 16639 22482 16677
rect 22282 16605 22298 16639
rect 22466 16605 22482 16639
rect 22282 16589 22482 16605
rect 22540 16639 22740 16677
rect 22798 16651 22998 16677
rect 23056 16651 23256 16677
rect 22540 16605 22556 16639
rect 22724 16605 22740 16639
rect 22540 16589 22740 16605
rect 23314 16639 23514 16677
rect 23314 16605 23330 16639
rect 23498 16605 23514 16639
rect 23314 16589 23514 16605
rect 23572 16639 23772 16677
rect 23572 16605 23588 16639
rect 23756 16605 23772 16639
rect 23572 16589 23772 16605
rect 20734 16513 20934 16529
rect 20734 16479 20750 16513
rect 20918 16479 20934 16513
rect 20734 16441 20934 16479
rect 20992 16513 21192 16529
rect 20992 16479 21008 16513
rect 21176 16479 21192 16513
rect 20992 16441 21192 16479
rect 21250 16513 21450 16529
rect 21250 16479 21266 16513
rect 21434 16479 21450 16513
rect 21250 16441 21450 16479
rect 21508 16513 21708 16529
rect 21508 16479 21524 16513
rect 21692 16479 21708 16513
rect 21508 16441 21708 16479
rect 21766 16513 21966 16529
rect 21766 16479 21782 16513
rect 21950 16479 21966 16513
rect 21766 16441 21966 16479
rect 22024 16513 22224 16529
rect 22024 16479 22040 16513
rect 22208 16479 22224 16513
rect 22024 16441 22224 16479
rect 22282 16513 22482 16529
rect 22282 16479 22298 16513
rect 22466 16479 22482 16513
rect 22282 16441 22482 16479
rect 22540 16513 22740 16529
rect 22540 16479 22556 16513
rect 22724 16479 22740 16513
rect 22540 16441 22740 16479
rect 22798 16513 22998 16529
rect 22798 16479 22814 16513
rect 22982 16479 22998 16513
rect 22798 16441 22998 16479
rect 23056 16513 23256 16529
rect 23056 16479 23072 16513
rect 23240 16479 23256 16513
rect 23056 16441 23256 16479
rect 23314 16513 23514 16529
rect 23314 16479 23330 16513
rect 23498 16479 23514 16513
rect 23314 16441 23514 16479
rect 23572 16513 23772 16529
rect 23572 16479 23588 16513
rect 23756 16479 23772 16513
rect 23572 16441 23772 16479
rect 20734 16331 20934 16357
rect 20992 16331 21192 16357
rect 21250 16331 21450 16357
rect 21508 16331 21708 16357
rect 21766 16331 21966 16357
rect 22024 16331 22224 16357
rect 22282 16331 22482 16357
rect 22540 16331 22740 16357
rect 22798 16331 22998 16357
rect 23056 16331 23256 16357
rect 23314 16331 23514 16357
rect 23572 16331 23772 16357
rect 12682 15407 12712 15429
rect 12766 15407 12796 15429
rect 12850 15407 12880 15429
rect 12934 15407 12964 15429
rect 13018 15407 13048 15429
rect 13102 15407 13132 15429
rect 13186 15407 13216 15429
rect 13270 15407 13300 15429
rect 12682 15251 12712 15277
rect 12766 15251 12796 15277
rect 12850 15251 12880 15277
rect 12934 15251 12964 15277
rect 13018 15251 13048 15277
rect 13102 15251 13132 15277
rect 13186 15251 13216 15277
rect 13270 15251 13300 15277
rect 26117 18009 26317 18035
rect 26375 18009 26575 18035
rect 26117 17771 26317 17809
rect 26117 17737 26133 17771
rect 26301 17737 26317 17771
rect 26117 17721 26317 17737
rect 26375 17771 26575 17809
rect 26375 17737 26391 17771
rect 26559 17737 26575 17771
rect 26375 17721 26575 17737
rect 26117 17126 26317 17142
rect 26117 17092 26133 17126
rect 26301 17092 26317 17126
rect 26117 17045 26317 17092
rect 26375 17126 26575 17142
rect 26375 17092 26391 17126
rect 26559 17092 26575 17126
rect 26375 17045 26575 17092
rect 26117 16819 26317 16845
rect 26375 16819 26575 16845
rect 26117 16549 26317 16575
rect 26375 16549 26575 16575
rect 26117 16311 26317 16349
rect 26117 16277 26133 16311
rect 26301 16277 26317 16311
rect 26117 16261 26317 16277
rect 26375 16311 26575 16349
rect 26375 16277 26391 16311
rect 26559 16277 26575 16311
rect 26375 16261 26575 16277
rect 25864 15597 25894 15623
rect 25948 15597 25978 15623
rect 26032 15597 26062 15623
rect 26116 15597 26146 15623
rect 26200 15597 26230 15623
rect 26284 15597 26314 15623
rect 26368 15597 26398 15623
rect 26452 15597 26482 15623
rect 25864 15365 25894 15397
rect 25948 15365 25978 15397
rect 26032 15365 26062 15397
rect 26116 15365 26146 15397
rect 26200 15365 26230 15397
rect 26284 15365 26314 15397
rect 26368 15365 26398 15397
rect 26452 15365 26482 15397
rect 25864 15349 26482 15365
rect 25864 15315 25904 15349
rect 25938 15315 25988 15349
rect 26022 15315 26072 15349
rect 26106 15315 26156 15349
rect 26190 15315 26240 15349
rect 26274 15315 26324 15349
rect 26358 15315 26408 15349
rect 26442 15315 26482 15349
rect 25864 15299 26482 15315
rect 25864 15277 25894 15299
rect 25948 15277 25978 15299
rect 26032 15277 26062 15299
rect 26116 15277 26146 15299
rect 26200 15277 26230 15299
rect 26284 15277 26314 15299
rect 26368 15277 26398 15299
rect 26452 15277 26482 15299
rect 25864 15121 25894 15147
rect 25948 15121 25978 15147
rect 26032 15121 26062 15147
rect 26116 15121 26146 15147
rect 26200 15121 26230 15147
rect 26284 15121 26314 15147
rect 26368 15121 26398 15147
rect 26452 15121 26482 15147
<< polycont >>
rect 12935 38358 13103 38392
rect 13193 38358 13361 38392
rect 25723 38476 25891 38510
rect 25981 38476 26149 38510
rect 7552 36829 7720 36863
rect 7810 36829 7978 36863
rect 8068 36829 8236 36863
rect 8326 36829 8494 36863
rect 8584 36829 8752 36863
rect 8842 36829 9010 36863
rect 9100 36829 9268 36863
rect 9358 36829 9526 36863
rect 9616 36829 9784 36863
rect 9874 36829 10042 36863
rect 10132 36829 10300 36863
rect 10390 36829 10558 36863
rect 7810 36721 7978 36755
rect 8584 36721 8752 36755
rect 8842 36721 9010 36755
rect 9616 36721 9784 36755
rect 9874 36721 10042 36755
rect 7552 36411 7720 36445
rect 8068 36411 8236 36445
rect 8326 36411 8494 36445
rect 9100 36411 9268 36445
rect 9358 36411 9526 36445
rect 10132 36411 10300 36445
rect 10390 36411 10558 36445
rect 7552 36285 7720 36319
rect 7810 36285 7978 36319
rect 8068 36285 8236 36319
rect 8326 36285 8494 36319
rect 8584 36285 8752 36319
rect 8842 36285 9010 36319
rect 9100 36285 9268 36319
rect 9358 36285 9526 36319
rect 9616 36285 9784 36319
rect 9874 36285 10042 36319
rect 10132 36285 10300 36319
rect 10390 36285 10558 36319
rect 12935 37543 13103 37577
rect 13193 37543 13361 37577
rect 12935 36898 13103 36932
rect 13193 36898 13361 36932
rect 12935 36083 13103 36117
rect 13193 36083 13361 36117
rect 20340 36947 20508 36981
rect 20598 36947 20766 36981
rect 20856 36947 21024 36981
rect 21114 36947 21282 36981
rect 21372 36947 21540 36981
rect 21630 36947 21798 36981
rect 21888 36947 22056 36981
rect 22146 36947 22314 36981
rect 22404 36947 22572 36981
rect 22662 36947 22830 36981
rect 22920 36947 23088 36981
rect 23178 36947 23346 36981
rect 20598 36839 20766 36873
rect 21372 36839 21540 36873
rect 21630 36839 21798 36873
rect 22404 36839 22572 36873
rect 22662 36839 22830 36873
rect 20340 36529 20508 36563
rect 20856 36529 21024 36563
rect 21114 36529 21282 36563
rect 21888 36529 22056 36563
rect 22146 36529 22314 36563
rect 22920 36529 23088 36563
rect 23178 36529 23346 36563
rect 20340 36403 20508 36437
rect 20598 36403 20766 36437
rect 20856 36403 21024 36437
rect 21114 36403 21282 36437
rect 21372 36403 21540 36437
rect 21630 36403 21798 36437
rect 21888 36403 22056 36437
rect 22146 36403 22314 36437
rect 22404 36403 22572 36437
rect 22662 36403 22830 36437
rect 22920 36403 23088 36437
rect 23178 36403 23346 36437
rect 12706 35121 12740 35155
rect 12790 35121 12824 35155
rect 12874 35121 12908 35155
rect 12958 35121 12992 35155
rect 13042 35121 13076 35155
rect 13126 35121 13160 35155
rect 13210 35121 13244 35155
rect 25723 37661 25891 37695
rect 25981 37661 26149 37695
rect 25723 37016 25891 37050
rect 25981 37016 26149 37050
rect 25723 36201 25891 36235
rect 25981 36201 26149 36235
rect 25494 35239 25528 35273
rect 25578 35239 25612 35273
rect 25662 35239 25696 35273
rect 25746 35239 25780 35273
rect 25830 35239 25864 35273
rect 25914 35239 25948 35273
rect 25998 35239 26032 35273
rect 12955 32432 13123 32466
rect 13213 32432 13381 32466
rect 25687 32356 25855 32390
rect 25945 32356 26113 32390
rect 7572 30903 7740 30937
rect 7830 30903 7998 30937
rect 8088 30903 8256 30937
rect 8346 30903 8514 30937
rect 8604 30903 8772 30937
rect 8862 30903 9030 30937
rect 9120 30903 9288 30937
rect 9378 30903 9546 30937
rect 9636 30903 9804 30937
rect 9894 30903 10062 30937
rect 10152 30903 10320 30937
rect 10410 30903 10578 30937
rect 7830 30795 7998 30829
rect 8604 30795 8772 30829
rect 8862 30795 9030 30829
rect 9636 30795 9804 30829
rect 9894 30795 10062 30829
rect 7572 30485 7740 30519
rect 8088 30485 8256 30519
rect 8346 30485 8514 30519
rect 9120 30485 9288 30519
rect 9378 30485 9546 30519
rect 10152 30485 10320 30519
rect 10410 30485 10578 30519
rect 7572 30359 7740 30393
rect 7830 30359 7998 30393
rect 8088 30359 8256 30393
rect 8346 30359 8514 30393
rect 8604 30359 8772 30393
rect 8862 30359 9030 30393
rect 9120 30359 9288 30393
rect 9378 30359 9546 30393
rect 9636 30359 9804 30393
rect 9894 30359 10062 30393
rect 10152 30359 10320 30393
rect 10410 30359 10578 30393
rect 12955 31617 13123 31651
rect 13213 31617 13381 31651
rect 12955 30972 13123 31006
rect 13213 30972 13381 31006
rect 12955 30157 13123 30191
rect 13213 30157 13381 30191
rect 20304 30827 20472 30861
rect 20562 30827 20730 30861
rect 20820 30827 20988 30861
rect 21078 30827 21246 30861
rect 21336 30827 21504 30861
rect 21594 30827 21762 30861
rect 21852 30827 22020 30861
rect 22110 30827 22278 30861
rect 22368 30827 22536 30861
rect 22626 30827 22794 30861
rect 22884 30827 23052 30861
rect 23142 30827 23310 30861
rect 20562 30719 20730 30753
rect 21336 30719 21504 30753
rect 21594 30719 21762 30753
rect 22368 30719 22536 30753
rect 22626 30719 22794 30753
rect 20304 30409 20472 30443
rect 20820 30409 20988 30443
rect 21078 30409 21246 30443
rect 21852 30409 22020 30443
rect 22110 30409 22278 30443
rect 22884 30409 23052 30443
rect 23142 30409 23310 30443
rect 20304 30283 20472 30317
rect 20562 30283 20730 30317
rect 20820 30283 20988 30317
rect 21078 30283 21246 30317
rect 21336 30283 21504 30317
rect 21594 30283 21762 30317
rect 21852 30283 22020 30317
rect 22110 30283 22278 30317
rect 22368 30283 22536 30317
rect 22626 30283 22794 30317
rect 22884 30283 23052 30317
rect 23142 30283 23310 30317
rect 12726 29195 12760 29229
rect 12810 29195 12844 29229
rect 12894 29195 12928 29229
rect 12978 29195 13012 29229
rect 13062 29195 13096 29229
rect 13146 29195 13180 29229
rect 13230 29195 13264 29229
rect 25687 31541 25855 31575
rect 25945 31541 26113 31575
rect 25687 30896 25855 30930
rect 25945 30896 26113 30930
rect 25687 30081 25855 30115
rect 25945 30081 26113 30115
rect 25458 29119 25492 29153
rect 25542 29119 25576 29153
rect 25626 29119 25660 29153
rect 25710 29119 25744 29153
rect 25794 29119 25828 29153
rect 25878 29119 25912 29153
rect 25962 29119 25996 29153
rect 13075 25728 13243 25762
rect 13333 25728 13501 25762
rect 25783 25598 25951 25632
rect 26041 25598 26209 25632
rect 7692 24199 7860 24233
rect 7950 24199 8118 24233
rect 8208 24199 8376 24233
rect 8466 24199 8634 24233
rect 8724 24199 8892 24233
rect 8982 24199 9150 24233
rect 9240 24199 9408 24233
rect 9498 24199 9666 24233
rect 9756 24199 9924 24233
rect 10014 24199 10182 24233
rect 10272 24199 10440 24233
rect 10530 24199 10698 24233
rect 7950 24091 8118 24125
rect 8724 24091 8892 24125
rect 8982 24091 9150 24125
rect 9756 24091 9924 24125
rect 10014 24091 10182 24125
rect 7692 23781 7860 23815
rect 8208 23781 8376 23815
rect 8466 23781 8634 23815
rect 9240 23781 9408 23815
rect 9498 23781 9666 23815
rect 10272 23781 10440 23815
rect 10530 23781 10698 23815
rect 7692 23655 7860 23689
rect 7950 23655 8118 23689
rect 8208 23655 8376 23689
rect 8466 23655 8634 23689
rect 8724 23655 8892 23689
rect 8982 23655 9150 23689
rect 9240 23655 9408 23689
rect 9498 23655 9666 23689
rect 9756 23655 9924 23689
rect 10014 23655 10182 23689
rect 10272 23655 10440 23689
rect 10530 23655 10698 23689
rect 13075 24913 13243 24947
rect 13333 24913 13501 24947
rect 13075 24268 13243 24302
rect 13333 24268 13501 24302
rect 13075 23453 13243 23487
rect 13333 23453 13501 23487
rect 12846 22491 12880 22525
rect 12930 22491 12964 22525
rect 13014 22491 13048 22525
rect 13098 22491 13132 22525
rect 13182 22491 13216 22525
rect 13266 22491 13300 22525
rect 13350 22491 13384 22525
rect 20400 24069 20568 24103
rect 20658 24069 20826 24103
rect 20916 24069 21084 24103
rect 21174 24069 21342 24103
rect 21432 24069 21600 24103
rect 21690 24069 21858 24103
rect 21948 24069 22116 24103
rect 22206 24069 22374 24103
rect 22464 24069 22632 24103
rect 22722 24069 22890 24103
rect 22980 24069 23148 24103
rect 23238 24069 23406 24103
rect 20658 23961 20826 23995
rect 21432 23961 21600 23995
rect 21690 23961 21858 23995
rect 22464 23961 22632 23995
rect 22722 23961 22890 23995
rect 20400 23651 20568 23685
rect 20916 23651 21084 23685
rect 21174 23651 21342 23685
rect 21948 23651 22116 23685
rect 22206 23651 22374 23685
rect 22980 23651 23148 23685
rect 23238 23651 23406 23685
rect 20400 23525 20568 23559
rect 20658 23525 20826 23559
rect 20916 23525 21084 23559
rect 21174 23525 21342 23559
rect 21432 23525 21600 23559
rect 21690 23525 21858 23559
rect 21948 23525 22116 23559
rect 22206 23525 22374 23559
rect 22464 23525 22632 23559
rect 22722 23525 22890 23559
rect 22980 23525 23148 23559
rect 23238 23525 23406 23559
rect 25783 24783 25951 24817
rect 26041 24783 26209 24817
rect 25783 24138 25951 24172
rect 26041 24138 26209 24172
rect 25783 23323 25951 23357
rect 26041 23323 26209 23357
rect 25554 22361 25588 22395
rect 25638 22361 25672 22395
rect 25722 22361 25756 22395
rect 25806 22361 25840 22395
rect 25890 22361 25924 22395
rect 25974 22361 26008 22395
rect 26058 22361 26092 22395
rect 12951 18682 13119 18716
rect 13209 18682 13377 18716
rect 26133 18552 26301 18586
rect 26391 18552 26559 18586
rect 7568 17153 7736 17187
rect 7826 17153 7994 17187
rect 8084 17153 8252 17187
rect 8342 17153 8510 17187
rect 8600 17153 8768 17187
rect 8858 17153 9026 17187
rect 9116 17153 9284 17187
rect 9374 17153 9542 17187
rect 9632 17153 9800 17187
rect 9890 17153 10058 17187
rect 10148 17153 10316 17187
rect 10406 17153 10574 17187
rect 7826 17045 7994 17079
rect 8600 17045 8768 17079
rect 8858 17045 9026 17079
rect 9632 17045 9800 17079
rect 9890 17045 10058 17079
rect 7568 16735 7736 16769
rect 8084 16735 8252 16769
rect 8342 16735 8510 16769
rect 9116 16735 9284 16769
rect 9374 16735 9542 16769
rect 10148 16735 10316 16769
rect 10406 16735 10574 16769
rect 7568 16609 7736 16643
rect 7826 16609 7994 16643
rect 8084 16609 8252 16643
rect 8342 16609 8510 16643
rect 8600 16609 8768 16643
rect 8858 16609 9026 16643
rect 9116 16609 9284 16643
rect 9374 16609 9542 16643
rect 9632 16609 9800 16643
rect 9890 16609 10058 16643
rect 10148 16609 10316 16643
rect 10406 16609 10574 16643
rect 12951 17867 13119 17901
rect 13209 17867 13377 17901
rect 12951 17222 13119 17256
rect 13209 17222 13377 17256
rect 12951 16407 13119 16441
rect 13209 16407 13377 16441
rect 12722 15445 12756 15479
rect 12806 15445 12840 15479
rect 12890 15445 12924 15479
rect 12974 15445 13008 15479
rect 13058 15445 13092 15479
rect 13142 15445 13176 15479
rect 13226 15445 13260 15479
rect 20750 17023 20918 17057
rect 21008 17023 21176 17057
rect 21266 17023 21434 17057
rect 21524 17023 21692 17057
rect 21782 17023 21950 17057
rect 22040 17023 22208 17057
rect 22298 17023 22466 17057
rect 22556 17023 22724 17057
rect 22814 17023 22982 17057
rect 23072 17023 23240 17057
rect 23330 17023 23498 17057
rect 23588 17023 23756 17057
rect 21008 16915 21176 16949
rect 21782 16915 21950 16949
rect 22040 16915 22208 16949
rect 22814 16915 22982 16949
rect 23072 16915 23240 16949
rect 20750 16605 20918 16639
rect 21266 16605 21434 16639
rect 21524 16605 21692 16639
rect 22298 16605 22466 16639
rect 22556 16605 22724 16639
rect 23330 16605 23498 16639
rect 23588 16605 23756 16639
rect 20750 16479 20918 16513
rect 21008 16479 21176 16513
rect 21266 16479 21434 16513
rect 21524 16479 21692 16513
rect 21782 16479 21950 16513
rect 22040 16479 22208 16513
rect 22298 16479 22466 16513
rect 22556 16479 22724 16513
rect 22814 16479 22982 16513
rect 23072 16479 23240 16513
rect 23330 16479 23498 16513
rect 23588 16479 23756 16513
rect 26133 17737 26301 17771
rect 26391 17737 26559 17771
rect 26133 17092 26301 17126
rect 26391 17092 26559 17126
rect 26133 16277 26301 16311
rect 26391 16277 26559 16311
rect 25904 15315 25938 15349
rect 25988 15315 26022 15349
rect 26072 15315 26106 15349
rect 26156 15315 26190 15349
rect 26240 15315 26274 15349
rect 26324 15315 26358 15349
rect 26408 15315 26442 15349
<< xpolycontact >>
rect 6892 37190 7324 37260
rect 6892 36028 7324 36098
rect 19680 37308 20112 37378
rect 19680 36146 20112 36216
rect 22410 34902 22842 35040
rect 23610 34902 24042 35040
rect 24410 37302 24548 37734
rect 24410 34902 24548 35334
rect 6912 31264 7344 31334
rect 6912 30102 7344 30172
rect 9642 28858 10074 28996
rect 10842 28858 11274 28996
rect 11642 31258 11780 31690
rect 11642 28858 11780 29290
rect 19644 31188 20076 31258
rect 19644 30026 20076 30096
rect 22374 28782 22806 28920
rect 23574 28782 24006 28920
rect 24374 31182 24512 31614
rect 24374 28782 24512 29214
rect 7032 24560 7464 24630
rect 7032 23398 7464 23468
rect 9762 22154 10194 22292
rect 10962 22154 11394 22292
rect 11762 24554 11900 24986
rect 11762 22154 11900 22586
rect 19740 24430 20172 24500
rect 19740 23268 20172 23338
rect 22470 22024 22902 22162
rect 23670 22024 24102 22162
rect 24470 24424 24608 24856
rect 24470 22024 24608 22456
rect 6908 17514 7340 17584
rect 6908 16352 7340 16422
rect 9638 15108 10070 15246
rect 10838 15108 11270 15246
rect 11638 17508 11776 17940
rect 11638 15108 11776 15540
rect 20090 17384 20522 17454
rect 20090 16222 20522 16292
rect 22820 14978 23252 15116
rect 24020 14978 24452 15116
rect 24820 17378 24958 17810
rect 24820 14978 24958 15410
<< xpolyres >>
rect 6188 37190 6892 37260
rect 6188 37094 6258 37190
rect 6188 37024 6788 37094
rect 6718 36928 6788 37024
rect 6188 36858 6788 36928
rect 6188 36762 6258 36858
rect 6188 36692 6788 36762
rect 6718 36596 6788 36692
rect 6188 36526 6788 36596
rect 6188 36430 6258 36526
rect 6188 36360 6788 36430
rect 6718 36264 6788 36360
rect 6188 36194 6788 36264
rect 6188 36098 6258 36194
rect 6188 36028 6892 36098
rect 18976 37308 19680 37378
rect 18976 37212 19046 37308
rect 18976 37142 19576 37212
rect 19506 37046 19576 37142
rect 18976 36976 19576 37046
rect 18976 36880 19046 36976
rect 18976 36810 19576 36880
rect 19506 36714 19576 36810
rect 18976 36644 19576 36714
rect 18976 36548 19046 36644
rect 18976 36478 19576 36548
rect 19506 36382 19576 36478
rect 18976 36312 19576 36382
rect 18976 36216 19046 36312
rect 18976 36146 19680 36216
rect 22842 34902 23610 35040
rect 24410 35334 24548 37302
rect 6208 31264 6912 31334
rect 6208 31168 6278 31264
rect 6208 31098 6808 31168
rect 6738 31002 6808 31098
rect 6208 30932 6808 31002
rect 6208 30836 6278 30932
rect 6208 30766 6808 30836
rect 6738 30670 6808 30766
rect 6208 30600 6808 30670
rect 6208 30504 6278 30600
rect 6208 30434 6808 30504
rect 6738 30338 6808 30434
rect 6208 30268 6808 30338
rect 6208 30172 6278 30268
rect 6208 30102 6912 30172
rect 10074 28858 10842 28996
rect 11642 29290 11780 31258
rect 18940 31188 19644 31258
rect 18940 31092 19010 31188
rect 18940 31022 19540 31092
rect 19470 30926 19540 31022
rect 18940 30856 19540 30926
rect 18940 30760 19010 30856
rect 18940 30690 19540 30760
rect 19470 30594 19540 30690
rect 18940 30524 19540 30594
rect 18940 30428 19010 30524
rect 18940 30358 19540 30428
rect 19470 30262 19540 30358
rect 18940 30192 19540 30262
rect 18940 30096 19010 30192
rect 18940 30026 19644 30096
rect 22806 28782 23574 28920
rect 24374 29214 24512 31182
rect 6328 24560 7032 24630
rect 6328 24464 6398 24560
rect 6328 24394 6928 24464
rect 6858 24298 6928 24394
rect 6328 24228 6928 24298
rect 6328 24132 6398 24228
rect 6328 24062 6928 24132
rect 6858 23966 6928 24062
rect 6328 23896 6928 23966
rect 6328 23800 6398 23896
rect 6328 23730 6928 23800
rect 6858 23634 6928 23730
rect 6328 23564 6928 23634
rect 6328 23468 6398 23564
rect 6328 23398 7032 23468
rect 10194 22154 10962 22292
rect 11762 22586 11900 24554
rect 19036 24430 19740 24500
rect 19036 24334 19106 24430
rect 19036 24264 19636 24334
rect 19566 24168 19636 24264
rect 19036 24098 19636 24168
rect 19036 24002 19106 24098
rect 19036 23932 19636 24002
rect 19566 23836 19636 23932
rect 19036 23766 19636 23836
rect 19036 23670 19106 23766
rect 19036 23600 19636 23670
rect 19566 23504 19636 23600
rect 19036 23434 19636 23504
rect 19036 23338 19106 23434
rect 19036 23268 19740 23338
rect 22902 22024 23670 22162
rect 24470 22456 24608 24424
rect 6204 17514 6908 17584
rect 6204 17418 6274 17514
rect 6204 17348 6804 17418
rect 6734 17252 6804 17348
rect 6204 17182 6804 17252
rect 6204 17086 6274 17182
rect 6204 17016 6804 17086
rect 6734 16920 6804 17016
rect 6204 16850 6804 16920
rect 6204 16754 6274 16850
rect 6204 16684 6804 16754
rect 6734 16588 6804 16684
rect 6204 16518 6804 16588
rect 6204 16422 6274 16518
rect 6204 16352 6908 16422
rect 10070 15108 10838 15246
rect 11638 15540 11776 17508
rect 19386 17384 20090 17454
rect 19386 17288 19456 17384
rect 19386 17218 19986 17288
rect 19916 17122 19986 17218
rect 19386 17052 19986 17122
rect 19386 16956 19456 17052
rect 19386 16886 19986 16956
rect 19916 16790 19986 16886
rect 19386 16720 19986 16790
rect 19386 16624 19456 16720
rect 19386 16554 19986 16624
rect 19916 16458 19986 16554
rect 19386 16388 19986 16458
rect 19386 16292 19456 16388
rect 19386 16222 20090 16292
rect 23252 14978 24020 15116
rect 24820 15410 24958 17378
<< locali >>
rect 25514 38613 26364 38626
rect 25514 38579 25643 38613
rect 26229 38579 26364 38613
rect 25514 38576 26364 38579
rect 25514 38516 25584 38576
rect 12726 38495 13576 38508
rect 12726 38461 12855 38495
rect 13441 38461 13576 38495
rect 12726 38458 13576 38461
rect 12726 38398 12796 38458
rect 12726 38096 12759 38398
rect 12793 38096 12796 38398
rect 13496 38398 13576 38458
rect 12919 38358 12935 38392
rect 13103 38358 13119 38392
rect 13177 38358 13193 38392
rect 13361 38358 13377 38392
rect 12873 38308 12907 38315
rect 12726 38058 12796 38096
rect 12856 38299 12926 38308
rect 12856 38123 12873 38299
rect 12907 38138 12926 38299
rect 13131 38299 13165 38315
rect 13389 38308 13423 38315
rect 12907 38123 13056 38138
rect 12856 38058 13056 38123
rect 13376 38299 13436 38308
rect 13376 38138 13389 38299
rect 13131 38107 13165 38123
rect 13236 38123 13389 38138
rect 13423 38123 13436 38299
rect 12996 37978 13056 38058
rect 13236 38058 13436 38123
rect 13496 38096 13503 38398
rect 13537 38338 13576 38398
rect 13537 38298 13776 38338
rect 13537 38118 13656 38298
rect 13756 38118 13776 38298
rect 25514 38214 25547 38516
rect 25581 38214 25584 38516
rect 26284 38516 26364 38576
rect 25707 38476 25723 38510
rect 25891 38476 25907 38510
rect 25965 38476 25981 38510
rect 26149 38476 26165 38510
rect 25661 38426 25695 38433
rect 25514 38176 25584 38214
rect 25644 38417 25714 38426
rect 25644 38241 25661 38417
rect 25695 38256 25714 38417
rect 25919 38417 25953 38433
rect 26177 38426 26211 38433
rect 25695 38241 25844 38256
rect 25644 38176 25844 38241
rect 26164 38417 26224 38426
rect 26164 38256 26177 38417
rect 25919 38225 25953 38241
rect 26024 38241 26177 38256
rect 26211 38241 26224 38417
rect 13537 38096 13776 38118
rect 13496 38078 13776 38096
rect 25784 38096 25844 38176
rect 26024 38176 26224 38241
rect 26284 38214 26291 38516
rect 26325 38456 26364 38516
rect 26325 38416 26564 38456
rect 26325 38236 26444 38416
rect 26544 38236 26564 38416
rect 26325 38214 26564 38236
rect 26284 38196 26564 38214
rect 26024 38096 26084 38176
rect 13236 37978 13296 38058
rect 5700 37938 11244 37948
rect 5700 35258 5716 37938
rect 5756 37882 11196 37898
rect 5756 35308 5766 37882
rect 5964 37608 10980 37618
rect 5964 35588 5976 37608
rect 6016 37552 10926 37568
rect 6016 35638 6030 37552
rect 6890 37260 10626 37278
rect 6890 37190 6892 37260
rect 7324 37238 10626 37260
rect 10576 37198 10626 37238
rect 7324 37190 10626 37198
rect 6890 37158 10626 37190
rect 7490 37098 7524 37114
rect 7490 36906 7524 36922
rect 7748 37098 7782 37114
rect 7748 36906 7782 36922
rect 8006 37098 8040 37114
rect 8006 36906 8040 36922
rect 8264 37098 8298 37114
rect 8264 36906 8298 36922
rect 8522 37098 8556 37114
rect 8522 36906 8556 36922
rect 8780 37098 8814 37114
rect 8780 36906 8814 36922
rect 9038 37098 9072 37114
rect 9038 36906 9072 36922
rect 9296 37098 9330 37114
rect 9296 36906 9330 36922
rect 9554 37098 9588 37114
rect 9554 36906 9588 36922
rect 9812 37098 9846 37114
rect 9812 36906 9846 36922
rect 10070 37098 10104 37114
rect 10070 36906 10104 36922
rect 10328 37098 10362 37114
rect 10328 36906 10362 36922
rect 10586 37098 10620 37114
rect 10586 36906 10620 36922
rect 7536 36829 7552 36863
rect 7720 36829 7736 36863
rect 7794 36829 7810 36863
rect 7978 36829 7994 36863
rect 8052 36829 8068 36863
rect 8236 36829 8252 36863
rect 8310 36829 8326 36863
rect 8494 36829 8510 36863
rect 8568 36829 8584 36863
rect 8752 36829 8768 36863
rect 8826 36829 8842 36863
rect 9010 36829 9026 36863
rect 9084 36829 9100 36863
rect 9268 36829 9284 36863
rect 9342 36829 9358 36863
rect 9526 36829 9542 36863
rect 9600 36829 9616 36863
rect 9784 36829 9800 36863
rect 9858 36829 9874 36863
rect 10042 36829 10058 36863
rect 10116 36829 10132 36863
rect 10300 36829 10316 36863
rect 10374 36829 10390 36863
rect 10558 36829 10574 36863
rect 7794 36721 7810 36755
rect 7978 36721 7994 36755
rect 8568 36721 8584 36755
rect 8752 36721 8768 36755
rect 8826 36721 8842 36755
rect 9010 36721 9026 36755
rect 9600 36721 9616 36755
rect 9784 36721 9800 36755
rect 9858 36721 9874 36755
rect 10042 36721 10058 36755
rect 7490 36671 7524 36687
rect 7490 36479 7524 36495
rect 7748 36671 7782 36687
rect 7748 36479 7782 36495
rect 8006 36671 8040 36687
rect 8006 36479 8040 36495
rect 8264 36671 8298 36687
rect 8264 36479 8298 36495
rect 8522 36671 8556 36687
rect 8522 36479 8556 36495
rect 8780 36671 8814 36687
rect 8780 36479 8814 36495
rect 9038 36671 9072 36687
rect 9038 36479 9072 36495
rect 9296 36671 9330 36687
rect 9296 36479 9330 36495
rect 9554 36671 9588 36687
rect 9554 36479 9588 36495
rect 9812 36671 9846 36687
rect 9812 36479 9846 36495
rect 10070 36671 10104 36687
rect 10070 36479 10104 36495
rect 10328 36671 10362 36687
rect 10328 36479 10362 36495
rect 10586 36671 10620 36687
rect 10586 36479 10620 36495
rect 7536 36411 7552 36445
rect 7720 36411 7736 36445
rect 8052 36411 8068 36445
rect 8236 36411 8252 36445
rect 8310 36411 8326 36445
rect 8494 36411 8510 36445
rect 9084 36411 9100 36445
rect 9268 36411 9284 36445
rect 9342 36411 9358 36445
rect 9526 36411 9542 36445
rect 10116 36411 10132 36445
rect 10300 36411 10316 36445
rect 10374 36411 10390 36445
rect 10558 36411 10574 36445
rect 7536 36285 7552 36319
rect 7720 36285 7736 36319
rect 7794 36285 7810 36319
rect 7978 36285 7994 36319
rect 8052 36285 8068 36319
rect 8236 36285 8252 36319
rect 8310 36285 8326 36319
rect 8494 36285 8510 36319
rect 8568 36285 8584 36319
rect 8752 36285 8768 36319
rect 8826 36285 8842 36319
rect 9010 36285 9026 36319
rect 9084 36285 9100 36319
rect 9268 36285 9284 36319
rect 9342 36285 9358 36319
rect 9526 36285 9542 36319
rect 9600 36285 9616 36319
rect 9784 36285 9800 36319
rect 9858 36285 9874 36319
rect 10042 36285 10058 36319
rect 10116 36285 10132 36319
rect 10300 36285 10316 36319
rect 10374 36285 10390 36319
rect 10558 36285 10574 36319
rect 7490 36235 7524 36251
rect 7490 36159 7524 36175
rect 7748 36235 7782 36251
rect 7748 36159 7782 36175
rect 8006 36235 8040 36251
rect 8006 36159 8040 36175
rect 8264 36235 8298 36251
rect 8264 36159 8298 36175
rect 8522 36235 8556 36251
rect 8522 36159 8556 36175
rect 8780 36235 8814 36251
rect 8780 36159 8814 36175
rect 9038 36235 9072 36251
rect 9038 36159 9072 36175
rect 9296 36235 9330 36251
rect 9296 36159 9330 36175
rect 9554 36235 9588 36251
rect 9554 36159 9588 36175
rect 9812 36235 9846 36251
rect 9812 36159 9846 36175
rect 10070 36235 10104 36251
rect 10070 36159 10104 36175
rect 10328 36235 10362 36251
rect 10328 36159 10362 36175
rect 10586 36235 10620 36251
rect 10586 36159 10620 36175
rect 6890 36108 7376 36138
rect 6890 36098 6956 36108
rect 6890 36028 6892 36098
rect 6890 36018 6956 36028
rect 7356 36018 7376 36108
rect 6890 35998 7376 36018
rect 7486 36048 10626 36078
rect 7486 35998 7526 36048
rect 10576 35998 10626 36048
rect 7486 35968 10626 35998
rect 10914 35638 10926 37552
rect 6016 35628 10926 35638
rect 10966 35588 10980 37608
rect 5964 35572 10980 35588
rect 11178 35308 11196 37882
rect 5756 35298 11196 35308
rect 11236 35258 11244 37938
rect 12996 37898 13296 37978
rect 18488 38056 24032 38066
rect 12726 37831 12796 37858
rect 11616 37598 11776 37618
rect 11616 37198 11636 37598
rect 11756 37198 11776 37598
rect 12726 37537 12759 37831
rect 12793 37537 12796 37831
rect 12856 37803 12926 37858
rect 12856 37658 12873 37803
rect 12907 37658 12926 37803
rect 13096 37803 13196 37898
rect 12873 37611 12907 37627
rect 13096 37627 13131 37803
rect 13165 37627 13196 37803
rect 13376 37803 13436 37858
rect 13376 37658 13389 37803
rect 13096 37618 13196 37627
rect 13423 37658 13436 37803
rect 13496 37831 13776 37858
rect 13131 37611 13165 37618
rect 13389 37611 13423 37627
rect 12919 37543 12935 37577
rect 13103 37543 13119 37577
rect 13177 37543 13193 37577
rect 13361 37543 13377 37577
rect 12726 37478 12796 37537
rect 13496 37537 13503 37831
rect 13537 37818 13776 37831
rect 13537 37638 13656 37818
rect 13756 37638 13776 37818
rect 13537 37598 13776 37638
rect 13537 37537 13576 37598
rect 13496 37478 13576 37537
rect 12726 37475 13576 37478
rect 12726 37441 12855 37475
rect 13441 37441 13576 37475
rect 12726 37408 13576 37441
rect 11616 37178 11776 37198
rect 12726 37035 13576 37048
rect 12726 37001 12855 37035
rect 13441 37001 13576 37035
rect 12726 36998 13576 37001
rect 12726 36938 12796 36998
rect 12726 36636 12759 36938
rect 12793 36636 12796 36938
rect 13496 36938 13576 36998
rect 12919 36898 12935 36932
rect 13103 36898 13119 36932
rect 13177 36898 13193 36932
rect 13361 36898 13377 36932
rect 12873 36848 12907 36855
rect 12726 36598 12796 36636
rect 12856 36839 12926 36848
rect 12856 36663 12873 36839
rect 12907 36678 12926 36839
rect 13131 36839 13165 36855
rect 13389 36848 13423 36855
rect 12907 36663 13056 36678
rect 12856 36598 13056 36663
rect 13376 36839 13436 36848
rect 13376 36678 13389 36839
rect 13131 36647 13165 36663
rect 13236 36663 13389 36678
rect 13423 36663 13436 36839
rect 12996 36518 13056 36598
rect 13236 36598 13436 36663
rect 13496 36636 13503 36938
rect 13537 36878 13576 36938
rect 13537 36838 13776 36878
rect 13537 36658 13656 36838
rect 13756 36658 13776 36838
rect 13537 36636 13776 36658
rect 13496 36618 13776 36636
rect 13236 36518 13296 36598
rect 12996 36438 13296 36518
rect 12726 36371 12796 36398
rect 12726 36077 12759 36371
rect 12793 36077 12796 36371
rect 12856 36343 12926 36398
rect 12856 36198 12873 36343
rect 12907 36198 12926 36343
rect 13096 36343 13196 36438
rect 12873 36151 12907 36167
rect 13096 36167 13131 36343
rect 13165 36167 13196 36343
rect 13376 36343 13436 36398
rect 13376 36198 13389 36343
rect 13096 36158 13196 36167
rect 13423 36198 13436 36343
rect 13496 36371 13776 36398
rect 13131 36151 13165 36158
rect 13389 36151 13423 36167
rect 12919 36083 12935 36117
rect 13103 36083 13119 36117
rect 13177 36083 13193 36117
rect 13361 36083 13377 36117
rect 12726 36018 12796 36077
rect 13496 36077 13503 36371
rect 13537 36358 13776 36371
rect 13537 36178 13656 36358
rect 13756 36178 13776 36358
rect 13537 36138 13776 36178
rect 13537 36077 13576 36138
rect 13496 36018 13576 36077
rect 12726 36015 13576 36018
rect 12726 35981 12855 36015
rect 13441 35981 13576 36015
rect 12726 35948 13576 35981
rect 12554 35433 12583 35467
rect 12617 35433 12675 35467
rect 12709 35433 12767 35467
rect 12801 35433 12859 35467
rect 12893 35433 12951 35467
rect 12985 35433 13043 35467
rect 13077 35433 13135 35467
rect 13169 35433 13227 35467
rect 13261 35433 13319 35467
rect 13353 35433 13411 35467
rect 13445 35433 13503 35467
rect 13537 35433 13566 35467
rect 12605 35391 12656 35433
rect 12605 35357 12622 35391
rect 12605 35323 12656 35357
rect 12605 35289 12622 35323
rect 12605 35273 12656 35289
rect 12690 35391 12756 35399
rect 12690 35357 12706 35391
rect 12740 35357 12756 35391
rect 12690 35323 12756 35357
rect 12690 35289 12706 35323
rect 12740 35289 12756 35323
rect 5700 35242 11244 35258
rect 12690 35255 12756 35289
rect 12790 35391 12824 35433
rect 12790 35323 12824 35357
rect 12790 35273 12824 35289
rect 12858 35391 12924 35399
rect 12858 35357 12874 35391
rect 12908 35357 12924 35391
rect 12858 35323 12924 35357
rect 12858 35289 12874 35323
rect 12908 35289 12924 35323
rect 12690 35239 12706 35255
rect 12571 35221 12706 35239
rect 12740 35239 12756 35255
rect 12858 35255 12924 35289
rect 12958 35391 12992 35433
rect 12958 35323 12992 35357
rect 12958 35273 12992 35289
rect 13026 35391 13092 35399
rect 13026 35357 13042 35391
rect 13076 35357 13092 35391
rect 13026 35323 13092 35357
rect 13026 35289 13042 35323
rect 13076 35289 13092 35323
rect 12858 35239 12874 35255
rect 12740 35221 12874 35239
rect 12908 35239 12924 35255
rect 13026 35255 13092 35289
rect 13126 35391 13160 35433
rect 13126 35323 13160 35357
rect 13126 35273 13160 35289
rect 13194 35391 13260 35399
rect 13194 35357 13210 35391
rect 13244 35357 13260 35391
rect 13194 35323 13260 35357
rect 13194 35289 13210 35323
rect 13244 35289 13260 35323
rect 13026 35239 13042 35255
rect 12908 35221 13042 35239
rect 13076 35239 13092 35255
rect 13194 35255 13260 35289
rect 13294 35391 13354 35433
rect 13328 35357 13354 35391
rect 13294 35323 13354 35357
rect 13328 35289 13354 35323
rect 13294 35273 13354 35289
rect 13399 35353 13549 35397
rect 18488 35376 18504 38056
rect 18544 38000 23984 38016
rect 18544 35426 18554 38000
rect 18752 37726 23768 37736
rect 18752 35706 18764 37726
rect 18804 37670 23714 37686
rect 18804 35756 18818 37670
rect 19678 37378 23414 37396
rect 19678 37308 19680 37378
rect 20112 37356 23414 37378
rect 23364 37316 23414 37356
rect 20112 37308 23414 37316
rect 19678 37276 23414 37308
rect 20278 37216 20312 37232
rect 20278 37024 20312 37040
rect 20536 37216 20570 37232
rect 20536 37024 20570 37040
rect 20794 37216 20828 37232
rect 20794 37024 20828 37040
rect 21052 37216 21086 37232
rect 21052 37024 21086 37040
rect 21310 37216 21344 37232
rect 21310 37024 21344 37040
rect 21568 37216 21602 37232
rect 21568 37024 21602 37040
rect 21826 37216 21860 37232
rect 21826 37024 21860 37040
rect 22084 37216 22118 37232
rect 22084 37024 22118 37040
rect 22342 37216 22376 37232
rect 22342 37024 22376 37040
rect 22600 37216 22634 37232
rect 22600 37024 22634 37040
rect 22858 37216 22892 37232
rect 22858 37024 22892 37040
rect 23116 37216 23150 37232
rect 23116 37024 23150 37040
rect 23374 37216 23408 37232
rect 23374 37024 23408 37040
rect 20324 36947 20340 36981
rect 20508 36947 20524 36981
rect 20582 36947 20598 36981
rect 20766 36947 20782 36981
rect 20840 36947 20856 36981
rect 21024 36947 21040 36981
rect 21098 36947 21114 36981
rect 21282 36947 21298 36981
rect 21356 36947 21372 36981
rect 21540 36947 21556 36981
rect 21614 36947 21630 36981
rect 21798 36947 21814 36981
rect 21872 36947 21888 36981
rect 22056 36947 22072 36981
rect 22130 36947 22146 36981
rect 22314 36947 22330 36981
rect 22388 36947 22404 36981
rect 22572 36947 22588 36981
rect 22646 36947 22662 36981
rect 22830 36947 22846 36981
rect 22904 36947 22920 36981
rect 23088 36947 23104 36981
rect 23162 36947 23178 36981
rect 23346 36947 23362 36981
rect 20582 36839 20598 36873
rect 20766 36839 20782 36873
rect 21356 36839 21372 36873
rect 21540 36839 21556 36873
rect 21614 36839 21630 36873
rect 21798 36839 21814 36873
rect 22388 36839 22404 36873
rect 22572 36839 22588 36873
rect 22646 36839 22662 36873
rect 22830 36839 22846 36873
rect 20278 36789 20312 36805
rect 20278 36597 20312 36613
rect 20536 36789 20570 36805
rect 20536 36597 20570 36613
rect 20794 36789 20828 36805
rect 20794 36597 20828 36613
rect 21052 36789 21086 36805
rect 21052 36597 21086 36613
rect 21310 36789 21344 36805
rect 21310 36597 21344 36613
rect 21568 36789 21602 36805
rect 21568 36597 21602 36613
rect 21826 36789 21860 36805
rect 21826 36597 21860 36613
rect 22084 36789 22118 36805
rect 22084 36597 22118 36613
rect 22342 36789 22376 36805
rect 22342 36597 22376 36613
rect 22600 36789 22634 36805
rect 22600 36597 22634 36613
rect 22858 36789 22892 36805
rect 22858 36597 22892 36613
rect 23116 36789 23150 36805
rect 23116 36597 23150 36613
rect 23374 36789 23408 36805
rect 23374 36597 23408 36613
rect 20324 36529 20340 36563
rect 20508 36529 20524 36563
rect 20840 36529 20856 36563
rect 21024 36529 21040 36563
rect 21098 36529 21114 36563
rect 21282 36529 21298 36563
rect 21872 36529 21888 36563
rect 22056 36529 22072 36563
rect 22130 36529 22146 36563
rect 22314 36529 22330 36563
rect 22904 36529 22920 36563
rect 23088 36529 23104 36563
rect 23162 36529 23178 36563
rect 23346 36529 23362 36563
rect 20324 36403 20340 36437
rect 20508 36403 20524 36437
rect 20582 36403 20598 36437
rect 20766 36403 20782 36437
rect 20840 36403 20856 36437
rect 21024 36403 21040 36437
rect 21098 36403 21114 36437
rect 21282 36403 21298 36437
rect 21356 36403 21372 36437
rect 21540 36403 21556 36437
rect 21614 36403 21630 36437
rect 21798 36403 21814 36437
rect 21872 36403 21888 36437
rect 22056 36403 22072 36437
rect 22130 36403 22146 36437
rect 22314 36403 22330 36437
rect 22388 36403 22404 36437
rect 22572 36403 22588 36437
rect 22646 36403 22662 36437
rect 22830 36403 22846 36437
rect 22904 36403 22920 36437
rect 23088 36403 23104 36437
rect 23162 36403 23178 36437
rect 23346 36403 23362 36437
rect 20278 36353 20312 36369
rect 20278 36277 20312 36293
rect 20536 36353 20570 36369
rect 20536 36277 20570 36293
rect 20794 36353 20828 36369
rect 20794 36277 20828 36293
rect 21052 36353 21086 36369
rect 21052 36277 21086 36293
rect 21310 36353 21344 36369
rect 21310 36277 21344 36293
rect 21568 36353 21602 36369
rect 21568 36277 21602 36293
rect 21826 36353 21860 36369
rect 21826 36277 21860 36293
rect 22084 36353 22118 36369
rect 22084 36277 22118 36293
rect 22342 36353 22376 36369
rect 22342 36277 22376 36293
rect 22600 36353 22634 36369
rect 22600 36277 22634 36293
rect 22858 36353 22892 36369
rect 22858 36277 22892 36293
rect 23116 36353 23150 36369
rect 23116 36277 23150 36293
rect 23374 36353 23408 36369
rect 23374 36277 23408 36293
rect 19678 36226 20164 36256
rect 19678 36216 19744 36226
rect 19678 36146 19680 36216
rect 19678 36136 19744 36146
rect 20144 36136 20164 36226
rect 19678 36116 20164 36136
rect 20274 36166 23414 36196
rect 20274 36116 20314 36166
rect 23364 36116 23414 36166
rect 20274 36086 23414 36116
rect 23702 35756 23714 37670
rect 18804 35746 23714 35756
rect 23754 35706 23768 37726
rect 18752 35690 23768 35706
rect 23966 35426 23984 38000
rect 18544 35416 23984 35426
rect 24024 35376 24032 38056
rect 25784 38016 26084 38096
rect 25514 37949 25584 37976
rect 24280 37830 24376 37864
rect 24582 37830 24678 37864
rect 24280 37768 24314 37830
rect 24204 36176 24280 36196
rect 24644 37768 24678 37830
rect 24404 37734 24564 37736
rect 24404 37302 24410 37734
rect 24548 37302 24564 37734
rect 24404 37296 24564 37302
rect 24314 36176 24344 36196
rect 24204 35736 24224 36176
rect 24324 35736 24344 36176
rect 24204 35716 24280 35736
rect 18488 35360 24032 35376
rect 13399 35319 13411 35353
rect 13445 35319 13503 35353
rect 13537 35319 13549 35353
rect 13194 35239 13210 35255
rect 13076 35221 13210 35239
rect 13244 35239 13260 35255
rect 13399 35269 13549 35319
rect 13244 35226 13365 35239
rect 13244 35221 13310 35226
rect 12571 35205 13310 35221
rect 12571 35087 12640 35205
rect 12690 35162 13261 35171
rect 12690 35128 12698 35162
rect 13186 35155 13261 35162
rect 13186 35128 13210 35155
rect 12690 35121 12706 35128
rect 12740 35121 12790 35128
rect 12824 35121 12874 35128
rect 12908 35121 12958 35128
rect 12992 35121 13042 35128
rect 13076 35121 13126 35128
rect 13160 35121 13210 35128
rect 13244 35121 13261 35155
rect 13301 35087 13310 35205
rect 12571 35067 13310 35087
rect 12571 35049 12706 35067
rect 12690 35033 12706 35049
rect 12740 35049 12874 35067
rect 12740 35033 12756 35049
rect 12605 34999 12656 35015
rect 12605 34965 12622 34999
rect 12605 34923 12656 34965
rect 12690 34999 12756 35033
rect 12858 35033 12874 35049
rect 12908 35049 13042 35067
rect 12908 35033 12924 35049
rect 12690 34965 12706 34999
rect 12740 34965 12756 34999
rect 12690 34957 12756 34965
rect 12790 34999 12824 35015
rect 12790 34923 12824 34965
rect 12858 34999 12924 35033
rect 13026 35033 13042 35049
rect 13076 35049 13210 35067
rect 13076 35033 13092 35049
rect 12858 34965 12874 34999
rect 12908 34965 12924 34999
rect 12858 34957 12924 34965
rect 12958 34999 12992 35015
rect 12958 34923 12992 34965
rect 13026 34999 13092 35033
rect 13194 35033 13210 35049
rect 13244 35062 13310 35067
rect 13358 35062 13365 35226
rect 13399 35235 13411 35269
rect 13445 35235 13503 35269
rect 13537 35235 13549 35269
rect 13399 35200 13549 35235
rect 22304 35176 23464 35196
rect 22304 35170 22324 35176
rect 23444 35170 23464 35176
rect 22280 35096 22324 35170
rect 24076 35136 24172 35170
rect 23444 35096 23464 35136
rect 22280 35076 23464 35096
rect 24138 35096 24172 35136
rect 22280 35074 22314 35076
rect 13244 35049 13365 35062
rect 13399 35051 13549 35068
rect 13244 35033 13260 35049
rect 13026 34965 13042 34999
rect 13076 34965 13092 34999
rect 13026 34957 13092 34965
rect 13126 34999 13160 35015
rect 13126 34923 13160 34965
rect 13194 34999 13260 35033
rect 13399 35017 13411 35051
rect 13445 35017 13503 35051
rect 13537 35017 13549 35051
rect 13194 34965 13210 34999
rect 13244 34965 13260 34999
rect 13194 34957 13260 34965
rect 13294 34999 13355 35015
rect 13328 34965 13355 34999
rect 13294 34923 13355 34965
rect 13399 34959 13549 35017
rect 12554 34889 12583 34923
rect 12617 34889 12675 34923
rect 12709 34889 12767 34923
rect 12801 34889 12859 34923
rect 12893 34889 12951 34923
rect 12985 34889 13043 34923
rect 13077 34889 13135 34923
rect 13169 34889 13227 34923
rect 13261 34889 13319 34923
rect 13353 34889 13411 34923
rect 13445 34889 13503 34923
rect 13537 34889 13566 34923
rect 24138 35074 24280 35096
rect 22280 34806 22314 34868
rect 24172 34868 24280 35074
rect 24314 35716 24344 35736
rect 24314 34868 24344 35096
rect 24138 34806 24344 34868
rect 25514 37655 25547 37949
rect 25581 37655 25584 37949
rect 25644 37921 25714 37976
rect 25644 37776 25661 37921
rect 25695 37776 25714 37921
rect 25884 37921 25984 38016
rect 25661 37729 25695 37745
rect 25884 37745 25919 37921
rect 25953 37745 25984 37921
rect 26164 37921 26224 37976
rect 26164 37776 26177 37921
rect 25884 37736 25984 37745
rect 26211 37776 26224 37921
rect 26284 37949 26564 37976
rect 25919 37729 25953 37736
rect 26177 37729 26211 37745
rect 25707 37661 25723 37695
rect 25891 37661 25907 37695
rect 25965 37661 25981 37695
rect 26149 37661 26165 37695
rect 25514 37596 25584 37655
rect 26284 37655 26291 37949
rect 26325 37936 26564 37949
rect 26325 37756 26444 37936
rect 26544 37756 26564 37936
rect 26325 37716 26564 37756
rect 26325 37655 26364 37716
rect 26284 37596 26364 37655
rect 25514 37593 26364 37596
rect 25514 37559 25643 37593
rect 26229 37559 26364 37593
rect 25514 37526 26364 37559
rect 25514 37153 26364 37166
rect 25514 37119 25643 37153
rect 26229 37119 26364 37153
rect 25514 37116 26364 37119
rect 25514 37056 25584 37116
rect 25514 36754 25547 37056
rect 25581 36754 25584 37056
rect 26284 37056 26364 37116
rect 25707 37016 25723 37050
rect 25891 37016 25907 37050
rect 25965 37016 25981 37050
rect 26149 37016 26165 37050
rect 25661 36966 25695 36973
rect 25514 36716 25584 36754
rect 25644 36957 25714 36966
rect 25644 36781 25661 36957
rect 25695 36796 25714 36957
rect 25919 36957 25953 36973
rect 26177 36966 26211 36973
rect 25695 36781 25844 36796
rect 25644 36716 25844 36781
rect 26164 36957 26224 36966
rect 26164 36796 26177 36957
rect 25919 36765 25953 36781
rect 26024 36781 26177 36796
rect 26211 36781 26224 36957
rect 25784 36636 25844 36716
rect 26024 36716 26224 36781
rect 26284 36754 26291 37056
rect 26325 36996 26364 37056
rect 26325 36956 26564 36996
rect 26325 36776 26444 36956
rect 26544 36776 26564 36956
rect 26325 36754 26564 36776
rect 26284 36736 26564 36754
rect 26024 36636 26084 36716
rect 25784 36556 26084 36636
rect 25514 36489 25584 36516
rect 25514 36195 25547 36489
rect 25581 36195 25584 36489
rect 25644 36461 25714 36516
rect 25644 36316 25661 36461
rect 25695 36316 25714 36461
rect 25884 36461 25984 36556
rect 25661 36269 25695 36285
rect 25884 36285 25919 36461
rect 25953 36285 25984 36461
rect 26164 36461 26224 36516
rect 26164 36316 26177 36461
rect 25884 36276 25984 36285
rect 26211 36316 26224 36461
rect 26284 36489 26564 36516
rect 25919 36269 25953 36276
rect 26177 36269 26211 36285
rect 25707 36201 25723 36235
rect 25891 36201 25907 36235
rect 25965 36201 25981 36235
rect 26149 36201 26165 36235
rect 25514 36136 25584 36195
rect 26284 36195 26291 36489
rect 26325 36476 26564 36489
rect 26325 36296 26444 36476
rect 26544 36296 26564 36476
rect 26325 36256 26564 36296
rect 26325 36195 26364 36256
rect 26284 36136 26364 36195
rect 25514 36133 26364 36136
rect 25514 36099 25643 36133
rect 26229 36099 26364 36133
rect 25514 36066 26364 36099
rect 25342 35551 25371 35585
rect 25405 35551 25463 35585
rect 25497 35551 25555 35585
rect 25589 35551 25647 35585
rect 25681 35551 25739 35585
rect 25773 35551 25831 35585
rect 25865 35551 25923 35585
rect 25957 35551 26015 35585
rect 26049 35551 26107 35585
rect 26141 35551 26199 35585
rect 26233 35551 26291 35585
rect 26325 35551 26354 35585
rect 25393 35509 25444 35551
rect 25393 35475 25410 35509
rect 25393 35441 25444 35475
rect 25393 35407 25410 35441
rect 25393 35391 25444 35407
rect 25478 35509 25544 35517
rect 25478 35475 25494 35509
rect 25528 35475 25544 35509
rect 25478 35441 25544 35475
rect 25478 35407 25494 35441
rect 25528 35407 25544 35441
rect 25478 35373 25544 35407
rect 25578 35509 25612 35551
rect 25578 35441 25612 35475
rect 25578 35391 25612 35407
rect 25646 35509 25712 35517
rect 25646 35475 25662 35509
rect 25696 35475 25712 35509
rect 25646 35441 25712 35475
rect 25646 35407 25662 35441
rect 25696 35407 25712 35441
rect 25478 35357 25494 35373
rect 25359 35339 25494 35357
rect 25528 35357 25544 35373
rect 25646 35373 25712 35407
rect 25746 35509 25780 35551
rect 25746 35441 25780 35475
rect 25746 35391 25780 35407
rect 25814 35509 25880 35517
rect 25814 35475 25830 35509
rect 25864 35475 25880 35509
rect 25814 35441 25880 35475
rect 25814 35407 25830 35441
rect 25864 35407 25880 35441
rect 25646 35357 25662 35373
rect 25528 35339 25662 35357
rect 25696 35357 25712 35373
rect 25814 35373 25880 35407
rect 25914 35509 25948 35551
rect 25914 35441 25948 35475
rect 25914 35391 25948 35407
rect 25982 35509 26048 35517
rect 25982 35475 25998 35509
rect 26032 35475 26048 35509
rect 25982 35441 26048 35475
rect 25982 35407 25998 35441
rect 26032 35407 26048 35441
rect 25814 35357 25830 35373
rect 25696 35339 25830 35357
rect 25864 35357 25880 35373
rect 25982 35373 26048 35407
rect 26082 35509 26142 35551
rect 26116 35475 26142 35509
rect 26082 35441 26142 35475
rect 26116 35407 26142 35441
rect 26082 35391 26142 35407
rect 26187 35471 26337 35515
rect 26187 35437 26199 35471
rect 26233 35437 26291 35471
rect 26325 35437 26337 35471
rect 25982 35357 25998 35373
rect 25864 35339 25998 35357
rect 26032 35357 26048 35373
rect 26187 35387 26337 35437
rect 26032 35344 26153 35357
rect 26032 35339 26098 35344
rect 25359 35323 26098 35339
rect 25359 35205 25428 35323
rect 25478 35280 26049 35289
rect 25478 35246 25486 35280
rect 25974 35273 26049 35280
rect 25974 35246 25998 35273
rect 25478 35239 25494 35246
rect 25528 35239 25578 35246
rect 25612 35239 25662 35246
rect 25696 35239 25746 35246
rect 25780 35239 25830 35246
rect 25864 35239 25914 35246
rect 25948 35239 25998 35246
rect 26032 35239 26049 35273
rect 26089 35205 26098 35323
rect 25359 35185 26098 35205
rect 25359 35167 25494 35185
rect 25478 35151 25494 35167
rect 25528 35167 25662 35185
rect 25528 35151 25544 35167
rect 25393 35117 25444 35133
rect 25393 35083 25410 35117
rect 25393 35041 25444 35083
rect 25478 35117 25544 35151
rect 25646 35151 25662 35167
rect 25696 35167 25830 35185
rect 25696 35151 25712 35167
rect 25478 35083 25494 35117
rect 25528 35083 25544 35117
rect 25478 35075 25544 35083
rect 25578 35117 25612 35133
rect 25578 35041 25612 35083
rect 25646 35117 25712 35151
rect 25814 35151 25830 35167
rect 25864 35167 25998 35185
rect 25864 35151 25880 35167
rect 25646 35083 25662 35117
rect 25696 35083 25712 35117
rect 25646 35075 25712 35083
rect 25746 35117 25780 35133
rect 25746 35041 25780 35083
rect 25814 35117 25880 35151
rect 25982 35151 25998 35167
rect 26032 35180 26098 35185
rect 26146 35180 26153 35344
rect 26187 35353 26199 35387
rect 26233 35353 26291 35387
rect 26325 35353 26337 35387
rect 26187 35318 26337 35353
rect 26032 35167 26153 35180
rect 26187 35169 26337 35186
rect 26032 35151 26048 35167
rect 25814 35083 25830 35117
rect 25864 35083 25880 35117
rect 25814 35075 25880 35083
rect 25914 35117 25948 35133
rect 25914 35041 25948 35083
rect 25982 35117 26048 35151
rect 26187 35135 26199 35169
rect 26233 35135 26291 35169
rect 26325 35135 26337 35169
rect 25982 35083 25998 35117
rect 26032 35083 26048 35117
rect 25982 35075 26048 35083
rect 26082 35117 26143 35133
rect 26116 35083 26143 35117
rect 26082 35041 26143 35083
rect 26187 35077 26337 35135
rect 25342 35007 25371 35041
rect 25405 35007 25463 35041
rect 25497 35007 25555 35041
rect 25589 35007 25647 35041
rect 25681 35007 25739 35041
rect 25773 35007 25831 35041
rect 25865 35007 25923 35041
rect 25957 35007 26015 35041
rect 26049 35007 26107 35041
rect 26141 35007 26199 35041
rect 26233 35007 26291 35041
rect 26325 35007 26354 35041
rect 24644 34806 24678 34868
rect 22280 34772 22376 34806
rect 24076 34776 24376 34806
rect 24076 34772 24172 34776
rect 24280 34772 24376 34776
rect 24582 34772 24678 34806
rect 12746 32569 13596 32582
rect 12746 32535 12875 32569
rect 13461 32535 13596 32569
rect 12746 32532 13596 32535
rect 12746 32472 12816 32532
rect 12746 32170 12779 32472
rect 12813 32170 12816 32472
rect 13516 32472 13596 32532
rect 12939 32432 12955 32466
rect 13123 32432 13139 32466
rect 13197 32432 13213 32466
rect 13381 32432 13397 32466
rect 12893 32382 12927 32389
rect 12746 32132 12816 32170
rect 12876 32373 12946 32382
rect 12876 32197 12893 32373
rect 12927 32212 12946 32373
rect 13151 32373 13185 32389
rect 13409 32382 13443 32389
rect 12927 32197 13076 32212
rect 12876 32132 13076 32197
rect 13396 32373 13456 32382
rect 13396 32212 13409 32373
rect 13151 32181 13185 32197
rect 13256 32197 13409 32212
rect 13443 32197 13456 32373
rect 13016 32052 13076 32132
rect 13256 32132 13456 32197
rect 13516 32170 13523 32472
rect 13557 32412 13596 32472
rect 25478 32493 26328 32506
rect 25478 32459 25607 32493
rect 26193 32459 26328 32493
rect 25478 32456 26328 32459
rect 13557 32372 13796 32412
rect 13557 32192 13676 32372
rect 13776 32192 13796 32372
rect 13557 32170 13796 32192
rect 13516 32152 13796 32170
rect 25478 32396 25548 32456
rect 13256 32052 13316 32132
rect 25478 32094 25511 32396
rect 25545 32094 25548 32396
rect 26248 32396 26328 32456
rect 25671 32356 25687 32390
rect 25855 32356 25871 32390
rect 25929 32356 25945 32390
rect 26113 32356 26129 32390
rect 25625 32306 25659 32313
rect 25478 32056 25548 32094
rect 25608 32297 25678 32306
rect 25608 32121 25625 32297
rect 25659 32136 25678 32297
rect 25883 32297 25917 32313
rect 26141 32306 26175 32313
rect 25659 32121 25808 32136
rect 25608 32056 25808 32121
rect 26128 32297 26188 32306
rect 26128 32136 26141 32297
rect 25883 32105 25917 32121
rect 25988 32121 26141 32136
rect 26175 32121 26188 32297
rect 5720 32012 11264 32022
rect 5720 29332 5736 32012
rect 5776 31956 11216 31972
rect 5776 29382 5786 31956
rect 5984 31682 11000 31692
rect 5984 29662 5996 31682
rect 6036 31626 10946 31642
rect 6036 29712 6050 31626
rect 6910 31334 10646 31352
rect 6910 31264 6912 31334
rect 7344 31312 10646 31334
rect 10596 31272 10646 31312
rect 7344 31264 10646 31272
rect 6910 31232 10646 31264
rect 7510 31172 7544 31188
rect 7510 30980 7544 30996
rect 7768 31172 7802 31188
rect 7768 30980 7802 30996
rect 8026 31172 8060 31188
rect 8026 30980 8060 30996
rect 8284 31172 8318 31188
rect 8284 30980 8318 30996
rect 8542 31172 8576 31188
rect 8542 30980 8576 30996
rect 8800 31172 8834 31188
rect 8800 30980 8834 30996
rect 9058 31172 9092 31188
rect 9058 30980 9092 30996
rect 9316 31172 9350 31188
rect 9316 30980 9350 30996
rect 9574 31172 9608 31188
rect 9574 30980 9608 30996
rect 9832 31172 9866 31188
rect 9832 30980 9866 30996
rect 10090 31172 10124 31188
rect 10090 30980 10124 30996
rect 10348 31172 10382 31188
rect 10348 30980 10382 30996
rect 10606 31172 10640 31188
rect 10606 30980 10640 30996
rect 7556 30903 7572 30937
rect 7740 30903 7756 30937
rect 7814 30903 7830 30937
rect 7998 30903 8014 30937
rect 8072 30903 8088 30937
rect 8256 30903 8272 30937
rect 8330 30903 8346 30937
rect 8514 30903 8530 30937
rect 8588 30903 8604 30937
rect 8772 30903 8788 30937
rect 8846 30903 8862 30937
rect 9030 30903 9046 30937
rect 9104 30903 9120 30937
rect 9288 30903 9304 30937
rect 9362 30903 9378 30937
rect 9546 30903 9562 30937
rect 9620 30903 9636 30937
rect 9804 30903 9820 30937
rect 9878 30903 9894 30937
rect 10062 30903 10078 30937
rect 10136 30903 10152 30937
rect 10320 30903 10336 30937
rect 10394 30903 10410 30937
rect 10578 30903 10594 30937
rect 7814 30795 7830 30829
rect 7998 30795 8014 30829
rect 8588 30795 8604 30829
rect 8772 30795 8788 30829
rect 8846 30795 8862 30829
rect 9030 30795 9046 30829
rect 9620 30795 9636 30829
rect 9804 30795 9820 30829
rect 9878 30795 9894 30829
rect 10062 30795 10078 30829
rect 7510 30745 7544 30761
rect 7510 30553 7544 30569
rect 7768 30745 7802 30761
rect 7768 30553 7802 30569
rect 8026 30745 8060 30761
rect 8026 30553 8060 30569
rect 8284 30745 8318 30761
rect 8284 30553 8318 30569
rect 8542 30745 8576 30761
rect 8542 30553 8576 30569
rect 8800 30745 8834 30761
rect 8800 30553 8834 30569
rect 9058 30745 9092 30761
rect 9058 30553 9092 30569
rect 9316 30745 9350 30761
rect 9316 30553 9350 30569
rect 9574 30745 9608 30761
rect 9574 30553 9608 30569
rect 9832 30745 9866 30761
rect 9832 30553 9866 30569
rect 10090 30745 10124 30761
rect 10090 30553 10124 30569
rect 10348 30745 10382 30761
rect 10348 30553 10382 30569
rect 10606 30745 10640 30761
rect 10606 30553 10640 30569
rect 7556 30485 7572 30519
rect 7740 30485 7756 30519
rect 8072 30485 8088 30519
rect 8256 30485 8272 30519
rect 8330 30485 8346 30519
rect 8514 30485 8530 30519
rect 9104 30485 9120 30519
rect 9288 30485 9304 30519
rect 9362 30485 9378 30519
rect 9546 30485 9562 30519
rect 10136 30485 10152 30519
rect 10320 30485 10336 30519
rect 10394 30485 10410 30519
rect 10578 30485 10594 30519
rect 7556 30359 7572 30393
rect 7740 30359 7756 30393
rect 7814 30359 7830 30393
rect 7998 30359 8014 30393
rect 8072 30359 8088 30393
rect 8256 30359 8272 30393
rect 8330 30359 8346 30393
rect 8514 30359 8530 30393
rect 8588 30359 8604 30393
rect 8772 30359 8788 30393
rect 8846 30359 8862 30393
rect 9030 30359 9046 30393
rect 9104 30359 9120 30393
rect 9288 30359 9304 30393
rect 9362 30359 9378 30393
rect 9546 30359 9562 30393
rect 9620 30359 9636 30393
rect 9804 30359 9820 30393
rect 9878 30359 9894 30393
rect 10062 30359 10078 30393
rect 10136 30359 10152 30393
rect 10320 30359 10336 30393
rect 10394 30359 10410 30393
rect 10578 30359 10594 30393
rect 7510 30309 7544 30325
rect 7510 30233 7544 30249
rect 7768 30309 7802 30325
rect 7768 30233 7802 30249
rect 8026 30309 8060 30325
rect 8026 30233 8060 30249
rect 8284 30309 8318 30325
rect 8284 30233 8318 30249
rect 8542 30309 8576 30325
rect 8542 30233 8576 30249
rect 8800 30309 8834 30325
rect 8800 30233 8834 30249
rect 9058 30309 9092 30325
rect 9058 30233 9092 30249
rect 9316 30309 9350 30325
rect 9316 30233 9350 30249
rect 9574 30309 9608 30325
rect 9574 30233 9608 30249
rect 9832 30309 9866 30325
rect 9832 30233 9866 30249
rect 10090 30309 10124 30325
rect 10090 30233 10124 30249
rect 10348 30309 10382 30325
rect 10348 30233 10382 30249
rect 10606 30309 10640 30325
rect 10606 30233 10640 30249
rect 6910 30182 7396 30212
rect 6910 30172 6976 30182
rect 6910 30102 6912 30172
rect 6910 30092 6976 30102
rect 7376 30092 7396 30182
rect 6910 30072 7396 30092
rect 7506 30122 10646 30152
rect 7506 30072 7546 30122
rect 10596 30072 10646 30122
rect 7506 30042 10646 30072
rect 10934 29712 10946 31626
rect 6036 29702 10946 29712
rect 10986 29662 11000 31682
rect 5984 29646 11000 29662
rect 11198 29382 11216 31956
rect 5776 29372 11216 29382
rect 11256 29332 11264 32012
rect 13016 31972 13316 32052
rect 25748 31976 25808 32056
rect 25988 32056 26188 32121
rect 26248 32094 26255 32396
rect 26289 32336 26328 32396
rect 26289 32296 26528 32336
rect 26289 32116 26408 32296
rect 26508 32116 26528 32296
rect 26289 32094 26528 32116
rect 26248 32076 26528 32094
rect 25988 31976 26048 32056
rect 12746 31905 12816 31932
rect 11512 31786 11608 31820
rect 11814 31786 11910 31820
rect 11512 31724 11546 31786
rect 11436 30132 11512 30152
rect 11876 31724 11910 31786
rect 11636 31690 11796 31692
rect 11636 31258 11642 31690
rect 11780 31258 11796 31690
rect 11636 31252 11796 31258
rect 11546 30132 11576 30152
rect 11436 29692 11456 30132
rect 11556 29692 11576 30132
rect 11436 29672 11512 29692
rect 5720 29316 11264 29332
rect 9536 29132 10696 29152
rect 9536 29126 9556 29132
rect 10676 29126 10696 29132
rect 9512 29052 9556 29126
rect 11308 29092 11404 29126
rect 10676 29052 10696 29092
rect 9512 29032 10696 29052
rect 11370 29052 11404 29092
rect 9512 29030 9546 29032
rect 11370 29030 11512 29052
rect 9512 28762 9546 28824
rect 11404 28824 11512 29030
rect 11546 29672 11576 29692
rect 11546 28824 11576 29052
rect 11370 28762 11576 28824
rect 12746 31611 12779 31905
rect 12813 31611 12816 31905
rect 12876 31877 12946 31932
rect 12876 31732 12893 31877
rect 12927 31732 12946 31877
rect 13116 31877 13216 31972
rect 18452 31936 23996 31946
rect 12893 31685 12927 31701
rect 13116 31701 13151 31877
rect 13185 31701 13216 31877
rect 13396 31877 13456 31932
rect 13396 31732 13409 31877
rect 13116 31692 13216 31701
rect 13443 31732 13456 31877
rect 13516 31905 13796 31932
rect 13151 31685 13185 31692
rect 13409 31685 13443 31701
rect 12939 31617 12955 31651
rect 13123 31617 13139 31651
rect 13197 31617 13213 31651
rect 13381 31617 13397 31651
rect 12746 31552 12816 31611
rect 13516 31611 13523 31905
rect 13557 31892 13796 31905
rect 13557 31712 13676 31892
rect 13776 31712 13796 31892
rect 13557 31672 13796 31712
rect 13557 31611 13596 31672
rect 13516 31552 13596 31611
rect 12746 31549 13596 31552
rect 12746 31515 12875 31549
rect 13461 31515 13596 31549
rect 12746 31482 13596 31515
rect 12746 31109 13596 31122
rect 12746 31075 12875 31109
rect 13461 31075 13596 31109
rect 12746 31072 13596 31075
rect 12746 31012 12816 31072
rect 12746 30710 12779 31012
rect 12813 30710 12816 31012
rect 13516 31012 13596 31072
rect 12939 30972 12955 31006
rect 13123 30972 13139 31006
rect 13197 30972 13213 31006
rect 13381 30972 13397 31006
rect 12893 30922 12927 30929
rect 12746 30672 12816 30710
rect 12876 30913 12946 30922
rect 12876 30737 12893 30913
rect 12927 30752 12946 30913
rect 13151 30913 13185 30929
rect 13409 30922 13443 30929
rect 12927 30737 13076 30752
rect 12876 30672 13076 30737
rect 13396 30913 13456 30922
rect 13396 30752 13409 30913
rect 13151 30721 13185 30737
rect 13256 30737 13409 30752
rect 13443 30737 13456 30913
rect 13016 30592 13076 30672
rect 13256 30672 13456 30737
rect 13516 30710 13523 31012
rect 13557 30952 13596 31012
rect 13557 30912 13796 30952
rect 13557 30732 13676 30912
rect 13776 30732 13796 30912
rect 13557 30710 13796 30732
rect 13516 30692 13796 30710
rect 13256 30592 13316 30672
rect 13016 30512 13316 30592
rect 12746 30445 12816 30472
rect 12746 30151 12779 30445
rect 12813 30151 12816 30445
rect 12876 30417 12946 30472
rect 12876 30272 12893 30417
rect 12927 30272 12946 30417
rect 13116 30417 13216 30512
rect 12893 30225 12927 30241
rect 13116 30241 13151 30417
rect 13185 30241 13216 30417
rect 13396 30417 13456 30472
rect 13396 30272 13409 30417
rect 13116 30232 13216 30241
rect 13443 30272 13456 30417
rect 13516 30445 13796 30472
rect 13151 30225 13185 30232
rect 13409 30225 13443 30241
rect 12939 30157 12955 30191
rect 13123 30157 13139 30191
rect 13197 30157 13213 30191
rect 13381 30157 13397 30191
rect 12746 30092 12816 30151
rect 13516 30151 13523 30445
rect 13557 30432 13796 30445
rect 13557 30252 13676 30432
rect 13776 30252 13796 30432
rect 13557 30212 13796 30252
rect 13557 30151 13596 30212
rect 13516 30092 13596 30151
rect 12746 30089 13596 30092
rect 12746 30055 12875 30089
rect 13461 30055 13596 30089
rect 12746 30022 13596 30055
rect 12574 29507 12603 29541
rect 12637 29507 12695 29541
rect 12729 29507 12787 29541
rect 12821 29507 12879 29541
rect 12913 29507 12971 29541
rect 13005 29507 13063 29541
rect 13097 29507 13155 29541
rect 13189 29507 13247 29541
rect 13281 29507 13339 29541
rect 13373 29507 13431 29541
rect 13465 29507 13523 29541
rect 13557 29507 13586 29541
rect 12625 29465 12676 29507
rect 12625 29431 12642 29465
rect 12625 29397 12676 29431
rect 12625 29363 12642 29397
rect 12625 29347 12676 29363
rect 12710 29465 12776 29473
rect 12710 29431 12726 29465
rect 12760 29431 12776 29465
rect 12710 29397 12776 29431
rect 12710 29363 12726 29397
rect 12760 29363 12776 29397
rect 12710 29329 12776 29363
rect 12810 29465 12844 29507
rect 12810 29397 12844 29431
rect 12810 29347 12844 29363
rect 12878 29465 12944 29473
rect 12878 29431 12894 29465
rect 12928 29431 12944 29465
rect 12878 29397 12944 29431
rect 12878 29363 12894 29397
rect 12928 29363 12944 29397
rect 12710 29313 12726 29329
rect 12591 29295 12726 29313
rect 12760 29313 12776 29329
rect 12878 29329 12944 29363
rect 12978 29465 13012 29507
rect 12978 29397 13012 29431
rect 12978 29347 13012 29363
rect 13046 29465 13112 29473
rect 13046 29431 13062 29465
rect 13096 29431 13112 29465
rect 13046 29397 13112 29431
rect 13046 29363 13062 29397
rect 13096 29363 13112 29397
rect 12878 29313 12894 29329
rect 12760 29295 12894 29313
rect 12928 29313 12944 29329
rect 13046 29329 13112 29363
rect 13146 29465 13180 29507
rect 13146 29397 13180 29431
rect 13146 29347 13180 29363
rect 13214 29465 13280 29473
rect 13214 29431 13230 29465
rect 13264 29431 13280 29465
rect 13214 29397 13280 29431
rect 13214 29363 13230 29397
rect 13264 29363 13280 29397
rect 13046 29313 13062 29329
rect 12928 29295 13062 29313
rect 13096 29313 13112 29329
rect 13214 29329 13280 29363
rect 13314 29465 13374 29507
rect 13348 29431 13374 29465
rect 13314 29397 13374 29431
rect 13348 29363 13374 29397
rect 13314 29347 13374 29363
rect 13419 29427 13569 29471
rect 13419 29393 13431 29427
rect 13465 29393 13523 29427
rect 13557 29393 13569 29427
rect 13214 29313 13230 29329
rect 13096 29295 13230 29313
rect 13264 29313 13280 29329
rect 13419 29343 13569 29393
rect 13264 29300 13385 29313
rect 13264 29295 13330 29300
rect 12591 29279 13330 29295
rect 12591 29161 12660 29279
rect 12710 29236 13281 29245
rect 12710 29202 12718 29236
rect 13206 29229 13281 29236
rect 13206 29202 13230 29229
rect 12710 29195 12726 29202
rect 12760 29195 12810 29202
rect 12844 29195 12894 29202
rect 12928 29195 12978 29202
rect 13012 29195 13062 29202
rect 13096 29195 13146 29202
rect 13180 29195 13230 29202
rect 13264 29195 13281 29229
rect 13321 29161 13330 29279
rect 12591 29141 13330 29161
rect 12591 29123 12726 29141
rect 12710 29107 12726 29123
rect 12760 29123 12894 29141
rect 12760 29107 12776 29123
rect 12625 29073 12676 29089
rect 12625 29039 12642 29073
rect 12625 28997 12676 29039
rect 12710 29073 12776 29107
rect 12878 29107 12894 29123
rect 12928 29123 13062 29141
rect 12928 29107 12944 29123
rect 12710 29039 12726 29073
rect 12760 29039 12776 29073
rect 12710 29031 12776 29039
rect 12810 29073 12844 29089
rect 12810 28997 12844 29039
rect 12878 29073 12944 29107
rect 13046 29107 13062 29123
rect 13096 29123 13230 29141
rect 13096 29107 13112 29123
rect 12878 29039 12894 29073
rect 12928 29039 12944 29073
rect 12878 29031 12944 29039
rect 12978 29073 13012 29089
rect 12978 28997 13012 29039
rect 13046 29073 13112 29107
rect 13214 29107 13230 29123
rect 13264 29136 13330 29141
rect 13378 29136 13385 29300
rect 13419 29309 13431 29343
rect 13465 29309 13523 29343
rect 13557 29309 13569 29343
rect 13419 29274 13569 29309
rect 18452 29256 18468 31936
rect 18508 31880 23948 31896
rect 18508 29306 18518 31880
rect 18716 31606 23732 31616
rect 18716 29586 18728 31606
rect 18768 31550 23678 31566
rect 18768 29636 18782 31550
rect 19642 31258 23378 31276
rect 19642 31188 19644 31258
rect 20076 31236 23378 31258
rect 23328 31196 23378 31236
rect 20076 31188 23378 31196
rect 19642 31156 23378 31188
rect 20242 31096 20276 31112
rect 20242 30904 20276 30920
rect 20500 31096 20534 31112
rect 20500 30904 20534 30920
rect 20758 31096 20792 31112
rect 20758 30904 20792 30920
rect 21016 31096 21050 31112
rect 21016 30904 21050 30920
rect 21274 31096 21308 31112
rect 21274 30904 21308 30920
rect 21532 31096 21566 31112
rect 21532 30904 21566 30920
rect 21790 31096 21824 31112
rect 21790 30904 21824 30920
rect 22048 31096 22082 31112
rect 22048 30904 22082 30920
rect 22306 31096 22340 31112
rect 22306 30904 22340 30920
rect 22564 31096 22598 31112
rect 22564 30904 22598 30920
rect 22822 31096 22856 31112
rect 22822 30904 22856 30920
rect 23080 31096 23114 31112
rect 23080 30904 23114 30920
rect 23338 31096 23372 31112
rect 23338 30904 23372 30920
rect 20288 30827 20304 30861
rect 20472 30827 20488 30861
rect 20546 30827 20562 30861
rect 20730 30827 20746 30861
rect 20804 30827 20820 30861
rect 20988 30827 21004 30861
rect 21062 30827 21078 30861
rect 21246 30827 21262 30861
rect 21320 30827 21336 30861
rect 21504 30827 21520 30861
rect 21578 30827 21594 30861
rect 21762 30827 21778 30861
rect 21836 30827 21852 30861
rect 22020 30827 22036 30861
rect 22094 30827 22110 30861
rect 22278 30827 22294 30861
rect 22352 30827 22368 30861
rect 22536 30827 22552 30861
rect 22610 30827 22626 30861
rect 22794 30827 22810 30861
rect 22868 30827 22884 30861
rect 23052 30827 23068 30861
rect 23126 30827 23142 30861
rect 23310 30827 23326 30861
rect 20546 30719 20562 30753
rect 20730 30719 20746 30753
rect 21320 30719 21336 30753
rect 21504 30719 21520 30753
rect 21578 30719 21594 30753
rect 21762 30719 21778 30753
rect 22352 30719 22368 30753
rect 22536 30719 22552 30753
rect 22610 30719 22626 30753
rect 22794 30719 22810 30753
rect 20242 30669 20276 30685
rect 20242 30477 20276 30493
rect 20500 30669 20534 30685
rect 20500 30477 20534 30493
rect 20758 30669 20792 30685
rect 20758 30477 20792 30493
rect 21016 30669 21050 30685
rect 21016 30477 21050 30493
rect 21274 30669 21308 30685
rect 21274 30477 21308 30493
rect 21532 30669 21566 30685
rect 21532 30477 21566 30493
rect 21790 30669 21824 30685
rect 21790 30477 21824 30493
rect 22048 30669 22082 30685
rect 22048 30477 22082 30493
rect 22306 30669 22340 30685
rect 22306 30477 22340 30493
rect 22564 30669 22598 30685
rect 22564 30477 22598 30493
rect 22822 30669 22856 30685
rect 22822 30477 22856 30493
rect 23080 30669 23114 30685
rect 23080 30477 23114 30493
rect 23338 30669 23372 30685
rect 23338 30477 23372 30493
rect 20288 30409 20304 30443
rect 20472 30409 20488 30443
rect 20804 30409 20820 30443
rect 20988 30409 21004 30443
rect 21062 30409 21078 30443
rect 21246 30409 21262 30443
rect 21836 30409 21852 30443
rect 22020 30409 22036 30443
rect 22094 30409 22110 30443
rect 22278 30409 22294 30443
rect 22868 30409 22884 30443
rect 23052 30409 23068 30443
rect 23126 30409 23142 30443
rect 23310 30409 23326 30443
rect 20288 30283 20304 30317
rect 20472 30283 20488 30317
rect 20546 30283 20562 30317
rect 20730 30283 20746 30317
rect 20804 30283 20820 30317
rect 20988 30283 21004 30317
rect 21062 30283 21078 30317
rect 21246 30283 21262 30317
rect 21320 30283 21336 30317
rect 21504 30283 21520 30317
rect 21578 30283 21594 30317
rect 21762 30283 21778 30317
rect 21836 30283 21852 30317
rect 22020 30283 22036 30317
rect 22094 30283 22110 30317
rect 22278 30283 22294 30317
rect 22352 30283 22368 30317
rect 22536 30283 22552 30317
rect 22610 30283 22626 30317
rect 22794 30283 22810 30317
rect 22868 30283 22884 30317
rect 23052 30283 23068 30317
rect 23126 30283 23142 30317
rect 23310 30283 23326 30317
rect 20242 30233 20276 30249
rect 20242 30157 20276 30173
rect 20500 30233 20534 30249
rect 20500 30157 20534 30173
rect 20758 30233 20792 30249
rect 20758 30157 20792 30173
rect 21016 30233 21050 30249
rect 21016 30157 21050 30173
rect 21274 30233 21308 30249
rect 21274 30157 21308 30173
rect 21532 30233 21566 30249
rect 21532 30157 21566 30173
rect 21790 30233 21824 30249
rect 21790 30157 21824 30173
rect 22048 30233 22082 30249
rect 22048 30157 22082 30173
rect 22306 30233 22340 30249
rect 22306 30157 22340 30173
rect 22564 30233 22598 30249
rect 22564 30157 22598 30173
rect 22822 30233 22856 30249
rect 22822 30157 22856 30173
rect 23080 30233 23114 30249
rect 23080 30157 23114 30173
rect 23338 30233 23372 30249
rect 23338 30157 23372 30173
rect 19642 30106 20128 30136
rect 19642 30096 19708 30106
rect 19642 30026 19644 30096
rect 19642 30016 19708 30026
rect 20108 30016 20128 30106
rect 19642 29996 20128 30016
rect 20238 30046 23378 30076
rect 20238 29996 20278 30046
rect 23328 29996 23378 30046
rect 20238 29966 23378 29996
rect 23666 29636 23678 31550
rect 18768 29626 23678 29636
rect 23718 29586 23732 31606
rect 18716 29570 23732 29586
rect 23930 29306 23948 31880
rect 18508 29296 23948 29306
rect 23988 29256 23996 31936
rect 25748 31896 26048 31976
rect 25478 31829 25548 31856
rect 24244 31710 24340 31744
rect 24546 31710 24642 31744
rect 24244 31648 24278 31710
rect 24168 30056 24244 30076
rect 24608 31648 24642 31710
rect 24368 31614 24528 31616
rect 24368 31182 24374 31614
rect 24512 31182 24528 31614
rect 24368 31176 24528 31182
rect 24278 30056 24308 30076
rect 24168 29616 24188 30056
rect 24288 29616 24308 30056
rect 24168 29596 24244 29616
rect 18452 29240 23996 29256
rect 13264 29123 13385 29136
rect 13419 29125 13569 29142
rect 13264 29107 13280 29123
rect 13046 29039 13062 29073
rect 13096 29039 13112 29073
rect 13046 29031 13112 29039
rect 13146 29073 13180 29089
rect 13146 28997 13180 29039
rect 13214 29073 13280 29107
rect 13419 29091 13431 29125
rect 13465 29091 13523 29125
rect 13557 29091 13569 29125
rect 13214 29039 13230 29073
rect 13264 29039 13280 29073
rect 13214 29031 13280 29039
rect 13314 29073 13375 29089
rect 13348 29039 13375 29073
rect 13314 28997 13375 29039
rect 13419 29033 13569 29091
rect 22268 29056 23428 29076
rect 22268 29050 22288 29056
rect 23408 29050 23428 29056
rect 12574 28963 12603 28997
rect 12637 28963 12695 28997
rect 12729 28963 12787 28997
rect 12821 28963 12879 28997
rect 12913 28963 12971 28997
rect 13005 28963 13063 28997
rect 13097 28963 13155 28997
rect 13189 28963 13247 28997
rect 13281 28963 13339 28997
rect 13373 28963 13431 28997
rect 13465 28963 13523 28997
rect 13557 28963 13586 28997
rect 22244 28976 22288 29050
rect 24040 29016 24136 29050
rect 23408 28976 23428 29016
rect 11876 28762 11910 28824
rect 9512 28728 9608 28762
rect 11308 28732 11608 28762
rect 11308 28728 11404 28732
rect 11512 28728 11608 28732
rect 11814 28728 11910 28762
rect 22244 28956 23428 28976
rect 24102 28976 24136 29016
rect 22244 28954 22278 28956
rect 24102 28954 24244 28976
rect 22244 28686 22278 28748
rect 24136 28748 24244 28954
rect 24278 29596 24308 29616
rect 24278 28748 24308 28976
rect 24102 28686 24308 28748
rect 25478 31535 25511 31829
rect 25545 31535 25548 31829
rect 25608 31801 25678 31856
rect 25608 31656 25625 31801
rect 25659 31656 25678 31801
rect 25848 31801 25948 31896
rect 25625 31609 25659 31625
rect 25848 31625 25883 31801
rect 25917 31625 25948 31801
rect 26128 31801 26188 31856
rect 26128 31656 26141 31801
rect 25848 31616 25948 31625
rect 26175 31656 26188 31801
rect 26248 31829 26528 31856
rect 25883 31609 25917 31616
rect 26141 31609 26175 31625
rect 25671 31541 25687 31575
rect 25855 31541 25871 31575
rect 25929 31541 25945 31575
rect 26113 31541 26129 31575
rect 25478 31476 25548 31535
rect 26248 31535 26255 31829
rect 26289 31816 26528 31829
rect 26289 31636 26408 31816
rect 26508 31636 26528 31816
rect 26289 31596 26528 31636
rect 26289 31535 26328 31596
rect 26248 31476 26328 31535
rect 25478 31473 26328 31476
rect 25478 31439 25607 31473
rect 26193 31439 26328 31473
rect 25478 31406 26328 31439
rect 25478 31033 26328 31046
rect 25478 30999 25607 31033
rect 26193 30999 26328 31033
rect 25478 30996 26328 30999
rect 25478 30936 25548 30996
rect 25478 30634 25511 30936
rect 25545 30634 25548 30936
rect 26248 30936 26328 30996
rect 25671 30896 25687 30930
rect 25855 30896 25871 30930
rect 25929 30896 25945 30930
rect 26113 30896 26129 30930
rect 25625 30846 25659 30853
rect 25478 30596 25548 30634
rect 25608 30837 25678 30846
rect 25608 30661 25625 30837
rect 25659 30676 25678 30837
rect 25883 30837 25917 30853
rect 26141 30846 26175 30853
rect 25659 30661 25808 30676
rect 25608 30596 25808 30661
rect 26128 30837 26188 30846
rect 26128 30676 26141 30837
rect 25883 30645 25917 30661
rect 25988 30661 26141 30676
rect 26175 30661 26188 30837
rect 25748 30516 25808 30596
rect 25988 30596 26188 30661
rect 26248 30634 26255 30936
rect 26289 30876 26328 30936
rect 26289 30836 26528 30876
rect 26289 30656 26408 30836
rect 26508 30656 26528 30836
rect 26289 30634 26528 30656
rect 26248 30616 26528 30634
rect 25988 30516 26048 30596
rect 25748 30436 26048 30516
rect 25478 30369 25548 30396
rect 25478 30075 25511 30369
rect 25545 30075 25548 30369
rect 25608 30341 25678 30396
rect 25608 30196 25625 30341
rect 25659 30196 25678 30341
rect 25848 30341 25948 30436
rect 25625 30149 25659 30165
rect 25848 30165 25883 30341
rect 25917 30165 25948 30341
rect 26128 30341 26188 30396
rect 26128 30196 26141 30341
rect 25848 30156 25948 30165
rect 26175 30196 26188 30341
rect 26248 30369 26528 30396
rect 25883 30149 25917 30156
rect 26141 30149 26175 30165
rect 25671 30081 25687 30115
rect 25855 30081 25871 30115
rect 25929 30081 25945 30115
rect 26113 30081 26129 30115
rect 25478 30016 25548 30075
rect 26248 30075 26255 30369
rect 26289 30356 26528 30369
rect 26289 30176 26408 30356
rect 26508 30176 26528 30356
rect 26289 30136 26528 30176
rect 26289 30075 26328 30136
rect 26248 30016 26328 30075
rect 25478 30013 26328 30016
rect 25478 29979 25607 30013
rect 26193 29979 26328 30013
rect 25478 29946 26328 29979
rect 25306 29431 25335 29465
rect 25369 29431 25427 29465
rect 25461 29431 25519 29465
rect 25553 29431 25611 29465
rect 25645 29431 25703 29465
rect 25737 29431 25795 29465
rect 25829 29431 25887 29465
rect 25921 29431 25979 29465
rect 26013 29431 26071 29465
rect 26105 29431 26163 29465
rect 26197 29431 26255 29465
rect 26289 29431 26318 29465
rect 25357 29389 25408 29431
rect 25357 29355 25374 29389
rect 25357 29321 25408 29355
rect 25357 29287 25374 29321
rect 25357 29271 25408 29287
rect 25442 29389 25508 29397
rect 25442 29355 25458 29389
rect 25492 29355 25508 29389
rect 25442 29321 25508 29355
rect 25442 29287 25458 29321
rect 25492 29287 25508 29321
rect 25442 29253 25508 29287
rect 25542 29389 25576 29431
rect 25542 29321 25576 29355
rect 25542 29271 25576 29287
rect 25610 29389 25676 29397
rect 25610 29355 25626 29389
rect 25660 29355 25676 29389
rect 25610 29321 25676 29355
rect 25610 29287 25626 29321
rect 25660 29287 25676 29321
rect 25442 29237 25458 29253
rect 25323 29219 25458 29237
rect 25492 29237 25508 29253
rect 25610 29253 25676 29287
rect 25710 29389 25744 29431
rect 25710 29321 25744 29355
rect 25710 29271 25744 29287
rect 25778 29389 25844 29397
rect 25778 29355 25794 29389
rect 25828 29355 25844 29389
rect 25778 29321 25844 29355
rect 25778 29287 25794 29321
rect 25828 29287 25844 29321
rect 25610 29237 25626 29253
rect 25492 29219 25626 29237
rect 25660 29237 25676 29253
rect 25778 29253 25844 29287
rect 25878 29389 25912 29431
rect 25878 29321 25912 29355
rect 25878 29271 25912 29287
rect 25946 29389 26012 29397
rect 25946 29355 25962 29389
rect 25996 29355 26012 29389
rect 25946 29321 26012 29355
rect 25946 29287 25962 29321
rect 25996 29287 26012 29321
rect 25778 29237 25794 29253
rect 25660 29219 25794 29237
rect 25828 29237 25844 29253
rect 25946 29253 26012 29287
rect 26046 29389 26106 29431
rect 26080 29355 26106 29389
rect 26046 29321 26106 29355
rect 26080 29287 26106 29321
rect 26046 29271 26106 29287
rect 26151 29351 26301 29395
rect 26151 29317 26163 29351
rect 26197 29317 26255 29351
rect 26289 29317 26301 29351
rect 25946 29237 25962 29253
rect 25828 29219 25962 29237
rect 25996 29237 26012 29253
rect 26151 29267 26301 29317
rect 25996 29224 26117 29237
rect 25996 29219 26062 29224
rect 25323 29203 26062 29219
rect 25323 29085 25392 29203
rect 25442 29160 26013 29169
rect 25442 29126 25450 29160
rect 25938 29153 26013 29160
rect 25938 29126 25962 29153
rect 25442 29119 25458 29126
rect 25492 29119 25542 29126
rect 25576 29119 25626 29126
rect 25660 29119 25710 29126
rect 25744 29119 25794 29126
rect 25828 29119 25878 29126
rect 25912 29119 25962 29126
rect 25996 29119 26013 29153
rect 26053 29085 26062 29203
rect 25323 29065 26062 29085
rect 25323 29047 25458 29065
rect 25442 29031 25458 29047
rect 25492 29047 25626 29065
rect 25492 29031 25508 29047
rect 25357 28997 25408 29013
rect 25357 28963 25374 28997
rect 25357 28921 25408 28963
rect 25442 28997 25508 29031
rect 25610 29031 25626 29047
rect 25660 29047 25794 29065
rect 25660 29031 25676 29047
rect 25442 28963 25458 28997
rect 25492 28963 25508 28997
rect 25442 28955 25508 28963
rect 25542 28997 25576 29013
rect 25542 28921 25576 28963
rect 25610 28997 25676 29031
rect 25778 29031 25794 29047
rect 25828 29047 25962 29065
rect 25828 29031 25844 29047
rect 25610 28963 25626 28997
rect 25660 28963 25676 28997
rect 25610 28955 25676 28963
rect 25710 28997 25744 29013
rect 25710 28921 25744 28963
rect 25778 28997 25844 29031
rect 25946 29031 25962 29047
rect 25996 29060 26062 29065
rect 26110 29060 26117 29224
rect 26151 29233 26163 29267
rect 26197 29233 26255 29267
rect 26289 29233 26301 29267
rect 26151 29198 26301 29233
rect 25996 29047 26117 29060
rect 26151 29049 26301 29066
rect 25996 29031 26012 29047
rect 25778 28963 25794 28997
rect 25828 28963 25844 28997
rect 25778 28955 25844 28963
rect 25878 28997 25912 29013
rect 25878 28921 25912 28963
rect 25946 28997 26012 29031
rect 26151 29015 26163 29049
rect 26197 29015 26255 29049
rect 26289 29015 26301 29049
rect 25946 28963 25962 28997
rect 25996 28963 26012 28997
rect 25946 28955 26012 28963
rect 26046 28997 26107 29013
rect 26080 28963 26107 28997
rect 26046 28921 26107 28963
rect 26151 28957 26301 29015
rect 25306 28887 25335 28921
rect 25369 28887 25427 28921
rect 25461 28887 25519 28921
rect 25553 28887 25611 28921
rect 25645 28887 25703 28921
rect 25737 28887 25795 28921
rect 25829 28887 25887 28921
rect 25921 28887 25979 28921
rect 26013 28887 26071 28921
rect 26105 28887 26163 28921
rect 26197 28887 26255 28921
rect 26289 28887 26318 28921
rect 24608 28686 24642 28748
rect 22244 28652 22340 28686
rect 24040 28656 24340 28686
rect 24040 28652 24136 28656
rect 24244 28652 24340 28656
rect 24546 28652 24642 28686
rect 12866 25865 13716 25878
rect 12866 25831 12995 25865
rect 13581 25831 13716 25865
rect 12866 25828 13716 25831
rect 12866 25768 12936 25828
rect 12866 25466 12899 25768
rect 12933 25466 12936 25768
rect 13636 25768 13716 25828
rect 13059 25728 13075 25762
rect 13243 25728 13259 25762
rect 13317 25728 13333 25762
rect 13501 25728 13517 25762
rect 13013 25678 13047 25685
rect 12866 25428 12936 25466
rect 12996 25669 13066 25678
rect 12996 25493 13013 25669
rect 13047 25508 13066 25669
rect 13271 25669 13305 25685
rect 13529 25678 13563 25685
rect 13047 25493 13196 25508
rect 12996 25428 13196 25493
rect 13516 25669 13576 25678
rect 13516 25508 13529 25669
rect 13271 25477 13305 25493
rect 13376 25493 13529 25508
rect 13563 25493 13576 25669
rect 13136 25348 13196 25428
rect 13376 25428 13576 25493
rect 13636 25466 13643 25768
rect 13677 25708 13716 25768
rect 25574 25735 26424 25748
rect 13677 25668 13916 25708
rect 13677 25488 13796 25668
rect 13896 25488 13916 25668
rect 13677 25466 13916 25488
rect 13636 25448 13916 25466
rect 25574 25701 25703 25735
rect 26289 25701 26424 25735
rect 25574 25698 26424 25701
rect 25574 25638 25644 25698
rect 13376 25348 13436 25428
rect 5840 25308 11384 25318
rect 5840 22628 5856 25308
rect 5896 25252 11336 25268
rect 5896 22678 5906 25252
rect 6104 24978 11120 24988
rect 6104 22958 6116 24978
rect 6156 24922 11066 24938
rect 6156 23008 6170 24922
rect 7030 24630 10766 24648
rect 7030 24560 7032 24630
rect 7464 24608 10766 24630
rect 10716 24568 10766 24608
rect 7464 24560 10766 24568
rect 7030 24528 10766 24560
rect 7630 24468 7664 24484
rect 7630 24276 7664 24292
rect 7888 24468 7922 24484
rect 7888 24276 7922 24292
rect 8146 24468 8180 24484
rect 8146 24276 8180 24292
rect 8404 24468 8438 24484
rect 8404 24276 8438 24292
rect 8662 24468 8696 24484
rect 8662 24276 8696 24292
rect 8920 24468 8954 24484
rect 8920 24276 8954 24292
rect 9178 24468 9212 24484
rect 9178 24276 9212 24292
rect 9436 24468 9470 24484
rect 9436 24276 9470 24292
rect 9694 24468 9728 24484
rect 9694 24276 9728 24292
rect 9952 24468 9986 24484
rect 9952 24276 9986 24292
rect 10210 24468 10244 24484
rect 10210 24276 10244 24292
rect 10468 24468 10502 24484
rect 10468 24276 10502 24292
rect 10726 24468 10760 24484
rect 10726 24276 10760 24292
rect 7676 24199 7692 24233
rect 7860 24199 7876 24233
rect 7934 24199 7950 24233
rect 8118 24199 8134 24233
rect 8192 24199 8208 24233
rect 8376 24199 8392 24233
rect 8450 24199 8466 24233
rect 8634 24199 8650 24233
rect 8708 24199 8724 24233
rect 8892 24199 8908 24233
rect 8966 24199 8982 24233
rect 9150 24199 9166 24233
rect 9224 24199 9240 24233
rect 9408 24199 9424 24233
rect 9482 24199 9498 24233
rect 9666 24199 9682 24233
rect 9740 24199 9756 24233
rect 9924 24199 9940 24233
rect 9998 24199 10014 24233
rect 10182 24199 10198 24233
rect 10256 24199 10272 24233
rect 10440 24199 10456 24233
rect 10514 24199 10530 24233
rect 10698 24199 10714 24233
rect 7934 24091 7950 24125
rect 8118 24091 8134 24125
rect 8708 24091 8724 24125
rect 8892 24091 8908 24125
rect 8966 24091 8982 24125
rect 9150 24091 9166 24125
rect 9740 24091 9756 24125
rect 9924 24091 9940 24125
rect 9998 24091 10014 24125
rect 10182 24091 10198 24125
rect 7630 24041 7664 24057
rect 7630 23849 7664 23865
rect 7888 24041 7922 24057
rect 7888 23849 7922 23865
rect 8146 24041 8180 24057
rect 8146 23849 8180 23865
rect 8404 24041 8438 24057
rect 8404 23849 8438 23865
rect 8662 24041 8696 24057
rect 8662 23849 8696 23865
rect 8920 24041 8954 24057
rect 8920 23849 8954 23865
rect 9178 24041 9212 24057
rect 9178 23849 9212 23865
rect 9436 24041 9470 24057
rect 9436 23849 9470 23865
rect 9694 24041 9728 24057
rect 9694 23849 9728 23865
rect 9952 24041 9986 24057
rect 9952 23849 9986 23865
rect 10210 24041 10244 24057
rect 10210 23849 10244 23865
rect 10468 24041 10502 24057
rect 10468 23849 10502 23865
rect 10726 24041 10760 24057
rect 10726 23849 10760 23865
rect 7676 23781 7692 23815
rect 7860 23781 7876 23815
rect 8192 23781 8208 23815
rect 8376 23781 8392 23815
rect 8450 23781 8466 23815
rect 8634 23781 8650 23815
rect 9224 23781 9240 23815
rect 9408 23781 9424 23815
rect 9482 23781 9498 23815
rect 9666 23781 9682 23815
rect 10256 23781 10272 23815
rect 10440 23781 10456 23815
rect 10514 23781 10530 23815
rect 10698 23781 10714 23815
rect 7676 23655 7692 23689
rect 7860 23655 7876 23689
rect 7934 23655 7950 23689
rect 8118 23655 8134 23689
rect 8192 23655 8208 23689
rect 8376 23655 8392 23689
rect 8450 23655 8466 23689
rect 8634 23655 8650 23689
rect 8708 23655 8724 23689
rect 8892 23655 8908 23689
rect 8966 23655 8982 23689
rect 9150 23655 9166 23689
rect 9224 23655 9240 23689
rect 9408 23655 9424 23689
rect 9482 23655 9498 23689
rect 9666 23655 9682 23689
rect 9740 23655 9756 23689
rect 9924 23655 9940 23689
rect 9998 23655 10014 23689
rect 10182 23655 10198 23689
rect 10256 23655 10272 23689
rect 10440 23655 10456 23689
rect 10514 23655 10530 23689
rect 10698 23655 10714 23689
rect 7630 23605 7664 23621
rect 7630 23529 7664 23545
rect 7888 23605 7922 23621
rect 7888 23529 7922 23545
rect 8146 23605 8180 23621
rect 8146 23529 8180 23545
rect 8404 23605 8438 23621
rect 8404 23529 8438 23545
rect 8662 23605 8696 23621
rect 8662 23529 8696 23545
rect 8920 23605 8954 23621
rect 8920 23529 8954 23545
rect 9178 23605 9212 23621
rect 9178 23529 9212 23545
rect 9436 23605 9470 23621
rect 9436 23529 9470 23545
rect 9694 23605 9728 23621
rect 9694 23529 9728 23545
rect 9952 23605 9986 23621
rect 9952 23529 9986 23545
rect 10210 23605 10244 23621
rect 10210 23529 10244 23545
rect 10468 23605 10502 23621
rect 10468 23529 10502 23545
rect 10726 23605 10760 23621
rect 10726 23529 10760 23545
rect 7030 23478 7516 23508
rect 7030 23468 7096 23478
rect 7030 23398 7032 23468
rect 7030 23388 7096 23398
rect 7496 23388 7516 23478
rect 7030 23368 7516 23388
rect 7626 23418 10766 23448
rect 7626 23368 7666 23418
rect 10716 23368 10766 23418
rect 7626 23338 10766 23368
rect 11054 23008 11066 24922
rect 6156 22998 11066 23008
rect 11106 22958 11120 24978
rect 6104 22942 11120 22958
rect 11318 22678 11336 25252
rect 5896 22668 11336 22678
rect 11376 22628 11384 25308
rect 13136 25268 13436 25348
rect 25574 25336 25607 25638
rect 25641 25336 25644 25638
rect 26344 25638 26424 25698
rect 25767 25598 25783 25632
rect 25951 25598 25967 25632
rect 26025 25598 26041 25632
rect 26209 25598 26225 25632
rect 25721 25548 25755 25555
rect 25574 25298 25644 25336
rect 25704 25539 25774 25548
rect 25704 25363 25721 25539
rect 25755 25378 25774 25539
rect 25979 25539 26013 25555
rect 26237 25548 26271 25555
rect 25755 25363 25904 25378
rect 25704 25298 25904 25363
rect 26224 25539 26284 25548
rect 26224 25378 26237 25539
rect 25979 25347 26013 25363
rect 26084 25363 26237 25378
rect 26271 25363 26284 25539
rect 12866 25201 12936 25228
rect 11632 25082 11728 25116
rect 11934 25082 12030 25116
rect 11632 25020 11666 25082
rect 11556 23428 11632 23448
rect 11996 25020 12030 25082
rect 11756 24986 11916 24988
rect 11756 24554 11762 24986
rect 11900 24554 11916 24986
rect 11756 24548 11916 24554
rect 11666 23428 11696 23448
rect 11556 22988 11576 23428
rect 11676 22988 11696 23428
rect 11556 22968 11632 22988
rect 5840 22612 11384 22628
rect 9656 22428 10816 22448
rect 9656 22422 9676 22428
rect 10796 22422 10816 22428
rect 9632 22348 9676 22422
rect 11428 22388 11524 22422
rect 10796 22348 10816 22388
rect 9632 22328 10816 22348
rect 11490 22348 11524 22388
rect 9632 22326 9666 22328
rect 11490 22326 11632 22348
rect 9632 22058 9666 22120
rect 11524 22120 11632 22326
rect 11666 22968 11696 22988
rect 11666 22120 11696 22348
rect 11490 22058 11696 22120
rect 12866 24907 12899 25201
rect 12933 24907 12936 25201
rect 12996 25173 13066 25228
rect 12996 25028 13013 25173
rect 13047 25028 13066 25173
rect 13236 25173 13336 25268
rect 13013 24981 13047 24997
rect 13236 24997 13271 25173
rect 13305 24997 13336 25173
rect 13516 25173 13576 25228
rect 13516 25028 13529 25173
rect 13236 24988 13336 24997
rect 13563 25028 13576 25173
rect 13636 25201 13916 25228
rect 13271 24981 13305 24988
rect 13529 24981 13563 24997
rect 13059 24913 13075 24947
rect 13243 24913 13259 24947
rect 13317 24913 13333 24947
rect 13501 24913 13517 24947
rect 12866 24848 12936 24907
rect 13636 24907 13643 25201
rect 13677 25188 13916 25201
rect 25844 25218 25904 25298
rect 26084 25298 26284 25363
rect 26344 25336 26351 25638
rect 26385 25578 26424 25638
rect 26385 25538 26624 25578
rect 26385 25358 26504 25538
rect 26604 25358 26624 25538
rect 26385 25336 26624 25358
rect 26344 25318 26624 25336
rect 26084 25218 26144 25298
rect 13677 25008 13796 25188
rect 13896 25008 13916 25188
rect 13677 24968 13916 25008
rect 18548 25178 24092 25188
rect 13677 24907 13716 24968
rect 13636 24848 13716 24907
rect 12866 24845 13716 24848
rect 12866 24811 12995 24845
rect 13581 24811 13716 24845
rect 12866 24778 13716 24811
rect 12866 24405 13716 24418
rect 12866 24371 12995 24405
rect 13581 24371 13716 24405
rect 12866 24368 13716 24371
rect 12866 24308 12936 24368
rect 12866 24006 12899 24308
rect 12933 24006 12936 24308
rect 13636 24308 13716 24368
rect 13059 24268 13075 24302
rect 13243 24268 13259 24302
rect 13317 24268 13333 24302
rect 13501 24268 13517 24302
rect 13013 24218 13047 24225
rect 12866 23968 12936 24006
rect 12996 24209 13066 24218
rect 12996 24033 13013 24209
rect 13047 24048 13066 24209
rect 13271 24209 13305 24225
rect 13529 24218 13563 24225
rect 13047 24033 13196 24048
rect 12996 23968 13196 24033
rect 13516 24209 13576 24218
rect 13516 24048 13529 24209
rect 13271 24017 13305 24033
rect 13376 24033 13529 24048
rect 13563 24033 13576 24209
rect 13136 23888 13196 23968
rect 13376 23968 13576 24033
rect 13636 24006 13643 24308
rect 13677 24248 13716 24308
rect 13677 24208 13916 24248
rect 13677 24028 13796 24208
rect 13896 24028 13916 24208
rect 13677 24006 13916 24028
rect 13636 23988 13916 24006
rect 13376 23888 13436 23968
rect 13136 23808 13436 23888
rect 12866 23741 12936 23768
rect 12866 23447 12899 23741
rect 12933 23447 12936 23741
rect 12996 23713 13066 23768
rect 12996 23568 13013 23713
rect 13047 23568 13066 23713
rect 13236 23713 13336 23808
rect 13013 23521 13047 23537
rect 13236 23537 13271 23713
rect 13305 23537 13336 23713
rect 13516 23713 13576 23768
rect 13516 23568 13529 23713
rect 13236 23528 13336 23537
rect 13563 23568 13576 23713
rect 13636 23741 13916 23768
rect 13271 23521 13305 23528
rect 13529 23521 13563 23537
rect 13059 23453 13075 23487
rect 13243 23453 13259 23487
rect 13317 23453 13333 23487
rect 13501 23453 13517 23487
rect 12866 23388 12936 23447
rect 13636 23447 13643 23741
rect 13677 23728 13916 23741
rect 13677 23548 13796 23728
rect 13896 23548 13916 23728
rect 13677 23508 13916 23548
rect 13677 23447 13716 23508
rect 13636 23388 13716 23447
rect 12866 23385 13716 23388
rect 12866 23351 12995 23385
rect 13581 23351 13716 23385
rect 12866 23318 13716 23351
rect 12694 22803 12723 22837
rect 12757 22803 12815 22837
rect 12849 22803 12907 22837
rect 12941 22803 12999 22837
rect 13033 22803 13091 22837
rect 13125 22803 13183 22837
rect 13217 22803 13275 22837
rect 13309 22803 13367 22837
rect 13401 22803 13459 22837
rect 13493 22803 13551 22837
rect 13585 22803 13643 22837
rect 13677 22803 13706 22837
rect 12745 22761 12796 22803
rect 12745 22727 12762 22761
rect 12745 22693 12796 22727
rect 12745 22659 12762 22693
rect 12745 22643 12796 22659
rect 12830 22761 12896 22769
rect 12830 22727 12846 22761
rect 12880 22727 12896 22761
rect 12830 22693 12896 22727
rect 12830 22659 12846 22693
rect 12880 22659 12896 22693
rect 12830 22625 12896 22659
rect 12930 22761 12964 22803
rect 12930 22693 12964 22727
rect 12930 22643 12964 22659
rect 12998 22761 13064 22769
rect 12998 22727 13014 22761
rect 13048 22727 13064 22761
rect 12998 22693 13064 22727
rect 12998 22659 13014 22693
rect 13048 22659 13064 22693
rect 12830 22609 12846 22625
rect 12711 22591 12846 22609
rect 12880 22609 12896 22625
rect 12998 22625 13064 22659
rect 13098 22761 13132 22803
rect 13098 22693 13132 22727
rect 13098 22643 13132 22659
rect 13166 22761 13232 22769
rect 13166 22727 13182 22761
rect 13216 22727 13232 22761
rect 13166 22693 13232 22727
rect 13166 22659 13182 22693
rect 13216 22659 13232 22693
rect 12998 22609 13014 22625
rect 12880 22591 13014 22609
rect 13048 22609 13064 22625
rect 13166 22625 13232 22659
rect 13266 22761 13300 22803
rect 13266 22693 13300 22727
rect 13266 22643 13300 22659
rect 13334 22761 13400 22769
rect 13334 22727 13350 22761
rect 13384 22727 13400 22761
rect 13334 22693 13400 22727
rect 13334 22659 13350 22693
rect 13384 22659 13400 22693
rect 13166 22609 13182 22625
rect 13048 22591 13182 22609
rect 13216 22609 13232 22625
rect 13334 22625 13400 22659
rect 13434 22761 13494 22803
rect 13468 22727 13494 22761
rect 13434 22693 13494 22727
rect 13468 22659 13494 22693
rect 13434 22643 13494 22659
rect 13539 22723 13689 22767
rect 13539 22689 13551 22723
rect 13585 22689 13643 22723
rect 13677 22689 13689 22723
rect 13334 22609 13350 22625
rect 13216 22591 13350 22609
rect 13384 22609 13400 22625
rect 13539 22639 13689 22689
rect 13384 22596 13505 22609
rect 13384 22591 13450 22596
rect 12711 22575 13450 22591
rect 12711 22457 12780 22575
rect 12830 22532 13401 22541
rect 12830 22498 12838 22532
rect 13326 22525 13401 22532
rect 13326 22498 13350 22525
rect 12830 22491 12846 22498
rect 12880 22491 12930 22498
rect 12964 22491 13014 22498
rect 13048 22491 13098 22498
rect 13132 22491 13182 22498
rect 13216 22491 13266 22498
rect 13300 22491 13350 22498
rect 13384 22491 13401 22525
rect 13441 22457 13450 22575
rect 12711 22437 13450 22457
rect 12711 22419 12846 22437
rect 12830 22403 12846 22419
rect 12880 22419 13014 22437
rect 12880 22403 12896 22419
rect 12745 22369 12796 22385
rect 12745 22335 12762 22369
rect 12745 22293 12796 22335
rect 12830 22369 12896 22403
rect 12998 22403 13014 22419
rect 13048 22419 13182 22437
rect 13048 22403 13064 22419
rect 12830 22335 12846 22369
rect 12880 22335 12896 22369
rect 12830 22327 12896 22335
rect 12930 22369 12964 22385
rect 12930 22293 12964 22335
rect 12998 22369 13064 22403
rect 13166 22403 13182 22419
rect 13216 22419 13350 22437
rect 13216 22403 13232 22419
rect 12998 22335 13014 22369
rect 13048 22335 13064 22369
rect 12998 22327 13064 22335
rect 13098 22369 13132 22385
rect 13098 22293 13132 22335
rect 13166 22369 13232 22403
rect 13334 22403 13350 22419
rect 13384 22432 13450 22437
rect 13498 22432 13505 22596
rect 13539 22605 13551 22639
rect 13585 22605 13643 22639
rect 13677 22605 13689 22639
rect 13539 22570 13689 22605
rect 18548 22498 18564 25178
rect 18604 25122 24044 25138
rect 18604 22548 18614 25122
rect 18812 24848 23828 24858
rect 18812 22828 18824 24848
rect 18864 24792 23774 24808
rect 18864 22878 18878 24792
rect 19738 24500 23474 24518
rect 19738 24430 19740 24500
rect 20172 24478 23474 24500
rect 23424 24438 23474 24478
rect 20172 24430 23474 24438
rect 19738 24398 23474 24430
rect 20338 24338 20372 24354
rect 20338 24146 20372 24162
rect 20596 24338 20630 24354
rect 20596 24146 20630 24162
rect 20854 24338 20888 24354
rect 20854 24146 20888 24162
rect 21112 24338 21146 24354
rect 21112 24146 21146 24162
rect 21370 24338 21404 24354
rect 21370 24146 21404 24162
rect 21628 24338 21662 24354
rect 21628 24146 21662 24162
rect 21886 24338 21920 24354
rect 21886 24146 21920 24162
rect 22144 24338 22178 24354
rect 22144 24146 22178 24162
rect 22402 24338 22436 24354
rect 22402 24146 22436 24162
rect 22660 24338 22694 24354
rect 22660 24146 22694 24162
rect 22918 24338 22952 24354
rect 22918 24146 22952 24162
rect 23176 24338 23210 24354
rect 23176 24146 23210 24162
rect 23434 24338 23468 24354
rect 23434 24146 23468 24162
rect 20384 24069 20400 24103
rect 20568 24069 20584 24103
rect 20642 24069 20658 24103
rect 20826 24069 20842 24103
rect 20900 24069 20916 24103
rect 21084 24069 21100 24103
rect 21158 24069 21174 24103
rect 21342 24069 21358 24103
rect 21416 24069 21432 24103
rect 21600 24069 21616 24103
rect 21674 24069 21690 24103
rect 21858 24069 21874 24103
rect 21932 24069 21948 24103
rect 22116 24069 22132 24103
rect 22190 24069 22206 24103
rect 22374 24069 22390 24103
rect 22448 24069 22464 24103
rect 22632 24069 22648 24103
rect 22706 24069 22722 24103
rect 22890 24069 22906 24103
rect 22964 24069 22980 24103
rect 23148 24069 23164 24103
rect 23222 24069 23238 24103
rect 23406 24069 23422 24103
rect 20642 23961 20658 23995
rect 20826 23961 20842 23995
rect 21416 23961 21432 23995
rect 21600 23961 21616 23995
rect 21674 23961 21690 23995
rect 21858 23961 21874 23995
rect 22448 23961 22464 23995
rect 22632 23961 22648 23995
rect 22706 23961 22722 23995
rect 22890 23961 22906 23995
rect 20338 23911 20372 23927
rect 20338 23719 20372 23735
rect 20596 23911 20630 23927
rect 20596 23719 20630 23735
rect 20854 23911 20888 23927
rect 20854 23719 20888 23735
rect 21112 23911 21146 23927
rect 21112 23719 21146 23735
rect 21370 23911 21404 23927
rect 21370 23719 21404 23735
rect 21628 23911 21662 23927
rect 21628 23719 21662 23735
rect 21886 23911 21920 23927
rect 21886 23719 21920 23735
rect 22144 23911 22178 23927
rect 22144 23719 22178 23735
rect 22402 23911 22436 23927
rect 22402 23719 22436 23735
rect 22660 23911 22694 23927
rect 22660 23719 22694 23735
rect 22918 23911 22952 23927
rect 22918 23719 22952 23735
rect 23176 23911 23210 23927
rect 23176 23719 23210 23735
rect 23434 23911 23468 23927
rect 23434 23719 23468 23735
rect 20384 23651 20400 23685
rect 20568 23651 20584 23685
rect 20900 23651 20916 23685
rect 21084 23651 21100 23685
rect 21158 23651 21174 23685
rect 21342 23651 21358 23685
rect 21932 23651 21948 23685
rect 22116 23651 22132 23685
rect 22190 23651 22206 23685
rect 22374 23651 22390 23685
rect 22964 23651 22980 23685
rect 23148 23651 23164 23685
rect 23222 23651 23238 23685
rect 23406 23651 23422 23685
rect 20384 23525 20400 23559
rect 20568 23525 20584 23559
rect 20642 23525 20658 23559
rect 20826 23525 20842 23559
rect 20900 23525 20916 23559
rect 21084 23525 21100 23559
rect 21158 23525 21174 23559
rect 21342 23525 21358 23559
rect 21416 23525 21432 23559
rect 21600 23525 21616 23559
rect 21674 23525 21690 23559
rect 21858 23525 21874 23559
rect 21932 23525 21948 23559
rect 22116 23525 22132 23559
rect 22190 23525 22206 23559
rect 22374 23525 22390 23559
rect 22448 23525 22464 23559
rect 22632 23525 22648 23559
rect 22706 23525 22722 23559
rect 22890 23525 22906 23559
rect 22964 23525 22980 23559
rect 23148 23525 23164 23559
rect 23222 23525 23238 23559
rect 23406 23525 23422 23559
rect 20338 23475 20372 23491
rect 20338 23399 20372 23415
rect 20596 23475 20630 23491
rect 20596 23399 20630 23415
rect 20854 23475 20888 23491
rect 20854 23399 20888 23415
rect 21112 23475 21146 23491
rect 21112 23399 21146 23415
rect 21370 23475 21404 23491
rect 21370 23399 21404 23415
rect 21628 23475 21662 23491
rect 21628 23399 21662 23415
rect 21886 23475 21920 23491
rect 21886 23399 21920 23415
rect 22144 23475 22178 23491
rect 22144 23399 22178 23415
rect 22402 23475 22436 23491
rect 22402 23399 22436 23415
rect 22660 23475 22694 23491
rect 22660 23399 22694 23415
rect 22918 23475 22952 23491
rect 22918 23399 22952 23415
rect 23176 23475 23210 23491
rect 23176 23399 23210 23415
rect 23434 23475 23468 23491
rect 23434 23399 23468 23415
rect 19738 23348 20224 23378
rect 19738 23338 19804 23348
rect 19738 23268 19740 23338
rect 19738 23258 19804 23268
rect 20204 23258 20224 23348
rect 19738 23238 20224 23258
rect 20334 23288 23474 23318
rect 20334 23238 20374 23288
rect 23424 23238 23474 23288
rect 20334 23208 23474 23238
rect 23762 22878 23774 24792
rect 18864 22868 23774 22878
rect 23814 22828 23828 24848
rect 18812 22812 23828 22828
rect 24026 22548 24044 25122
rect 18604 22538 24044 22548
rect 24084 22498 24092 25178
rect 25844 25138 26144 25218
rect 25574 25071 25644 25098
rect 24340 24952 24436 24986
rect 24642 24952 24738 24986
rect 24340 24890 24374 24952
rect 24264 23298 24340 23318
rect 24704 24890 24738 24952
rect 24464 24856 24624 24858
rect 24464 24424 24470 24856
rect 24608 24424 24624 24856
rect 24464 24418 24624 24424
rect 24374 23298 24404 23318
rect 24264 22858 24284 23298
rect 24384 22858 24404 23298
rect 24264 22838 24340 22858
rect 18548 22482 24092 22498
rect 13384 22419 13505 22432
rect 13539 22421 13689 22438
rect 13384 22403 13400 22419
rect 13166 22335 13182 22369
rect 13216 22335 13232 22369
rect 13166 22327 13232 22335
rect 13266 22369 13300 22385
rect 13266 22293 13300 22335
rect 13334 22369 13400 22403
rect 13539 22387 13551 22421
rect 13585 22387 13643 22421
rect 13677 22387 13689 22421
rect 13334 22335 13350 22369
rect 13384 22335 13400 22369
rect 13334 22327 13400 22335
rect 13434 22369 13495 22385
rect 13468 22335 13495 22369
rect 13434 22293 13495 22335
rect 13539 22329 13689 22387
rect 22364 22298 23524 22318
rect 12694 22259 12723 22293
rect 12757 22259 12815 22293
rect 12849 22259 12907 22293
rect 12941 22259 12999 22293
rect 13033 22259 13091 22293
rect 13125 22259 13183 22293
rect 13217 22259 13275 22293
rect 13309 22259 13367 22293
rect 13401 22259 13459 22293
rect 13493 22259 13551 22293
rect 13585 22259 13643 22293
rect 13677 22259 13706 22293
rect 22364 22292 22384 22298
rect 23504 22292 23524 22298
rect 11996 22058 12030 22120
rect 9632 22024 9728 22058
rect 11428 22028 11728 22058
rect 11428 22024 11524 22028
rect 11632 22024 11728 22028
rect 11934 22024 12030 22058
rect 22340 22218 22384 22292
rect 24136 22258 24232 22292
rect 23504 22218 23524 22258
rect 22340 22198 23524 22218
rect 24198 22218 24232 22258
rect 22340 22196 22374 22198
rect 24198 22196 24340 22218
rect 22340 21928 22374 21990
rect 24232 21990 24340 22196
rect 24374 22838 24404 22858
rect 24374 21990 24404 22218
rect 24198 21928 24404 21990
rect 25574 24777 25607 25071
rect 25641 24777 25644 25071
rect 25704 25043 25774 25098
rect 25704 24898 25721 25043
rect 25755 24898 25774 25043
rect 25944 25043 26044 25138
rect 25721 24851 25755 24867
rect 25944 24867 25979 25043
rect 26013 24867 26044 25043
rect 26224 25043 26284 25098
rect 26224 24898 26237 25043
rect 25944 24858 26044 24867
rect 26271 24898 26284 25043
rect 26344 25071 26624 25098
rect 25979 24851 26013 24858
rect 26237 24851 26271 24867
rect 25767 24783 25783 24817
rect 25951 24783 25967 24817
rect 26025 24783 26041 24817
rect 26209 24783 26225 24817
rect 25574 24718 25644 24777
rect 26344 24777 26351 25071
rect 26385 25058 26624 25071
rect 26385 24878 26504 25058
rect 26604 24878 26624 25058
rect 26385 24838 26624 24878
rect 26385 24777 26424 24838
rect 26344 24718 26424 24777
rect 25574 24715 26424 24718
rect 25574 24681 25703 24715
rect 26289 24681 26424 24715
rect 25574 24648 26424 24681
rect 25574 24275 26424 24288
rect 25574 24241 25703 24275
rect 26289 24241 26424 24275
rect 25574 24238 26424 24241
rect 25574 24178 25644 24238
rect 25574 23876 25607 24178
rect 25641 23876 25644 24178
rect 26344 24178 26424 24238
rect 25767 24138 25783 24172
rect 25951 24138 25967 24172
rect 26025 24138 26041 24172
rect 26209 24138 26225 24172
rect 25721 24088 25755 24095
rect 25574 23838 25644 23876
rect 25704 24079 25774 24088
rect 25704 23903 25721 24079
rect 25755 23918 25774 24079
rect 25979 24079 26013 24095
rect 26237 24088 26271 24095
rect 25755 23903 25904 23918
rect 25704 23838 25904 23903
rect 26224 24079 26284 24088
rect 26224 23918 26237 24079
rect 25979 23887 26013 23903
rect 26084 23903 26237 23918
rect 26271 23903 26284 24079
rect 25844 23758 25904 23838
rect 26084 23838 26284 23903
rect 26344 23876 26351 24178
rect 26385 24118 26424 24178
rect 26385 24078 26624 24118
rect 26385 23898 26504 24078
rect 26604 23898 26624 24078
rect 26385 23876 26624 23898
rect 26344 23858 26624 23876
rect 26084 23758 26144 23838
rect 25844 23678 26144 23758
rect 25574 23611 25644 23638
rect 25574 23317 25607 23611
rect 25641 23317 25644 23611
rect 25704 23583 25774 23638
rect 25704 23438 25721 23583
rect 25755 23438 25774 23583
rect 25944 23583 26044 23678
rect 25721 23391 25755 23407
rect 25944 23407 25979 23583
rect 26013 23407 26044 23583
rect 26224 23583 26284 23638
rect 26224 23438 26237 23583
rect 25944 23398 26044 23407
rect 26271 23438 26284 23583
rect 26344 23611 26624 23638
rect 25979 23391 26013 23398
rect 26237 23391 26271 23407
rect 25767 23323 25783 23357
rect 25951 23323 25967 23357
rect 26025 23323 26041 23357
rect 26209 23323 26225 23357
rect 25574 23258 25644 23317
rect 26344 23317 26351 23611
rect 26385 23598 26624 23611
rect 26385 23418 26504 23598
rect 26604 23418 26624 23598
rect 26385 23378 26624 23418
rect 26385 23317 26424 23378
rect 26344 23258 26424 23317
rect 25574 23255 26424 23258
rect 25574 23221 25703 23255
rect 26289 23221 26424 23255
rect 25574 23188 26424 23221
rect 25402 22673 25431 22707
rect 25465 22673 25523 22707
rect 25557 22673 25615 22707
rect 25649 22673 25707 22707
rect 25741 22673 25799 22707
rect 25833 22673 25891 22707
rect 25925 22673 25983 22707
rect 26017 22673 26075 22707
rect 26109 22673 26167 22707
rect 26201 22673 26259 22707
rect 26293 22673 26351 22707
rect 26385 22673 26414 22707
rect 25453 22631 25504 22673
rect 25453 22597 25470 22631
rect 25453 22563 25504 22597
rect 25453 22529 25470 22563
rect 25453 22513 25504 22529
rect 25538 22631 25604 22639
rect 25538 22597 25554 22631
rect 25588 22597 25604 22631
rect 25538 22563 25604 22597
rect 25538 22529 25554 22563
rect 25588 22529 25604 22563
rect 25538 22495 25604 22529
rect 25638 22631 25672 22673
rect 25638 22563 25672 22597
rect 25638 22513 25672 22529
rect 25706 22631 25772 22639
rect 25706 22597 25722 22631
rect 25756 22597 25772 22631
rect 25706 22563 25772 22597
rect 25706 22529 25722 22563
rect 25756 22529 25772 22563
rect 25538 22479 25554 22495
rect 25419 22461 25554 22479
rect 25588 22479 25604 22495
rect 25706 22495 25772 22529
rect 25806 22631 25840 22673
rect 25806 22563 25840 22597
rect 25806 22513 25840 22529
rect 25874 22631 25940 22639
rect 25874 22597 25890 22631
rect 25924 22597 25940 22631
rect 25874 22563 25940 22597
rect 25874 22529 25890 22563
rect 25924 22529 25940 22563
rect 25706 22479 25722 22495
rect 25588 22461 25722 22479
rect 25756 22479 25772 22495
rect 25874 22495 25940 22529
rect 25974 22631 26008 22673
rect 25974 22563 26008 22597
rect 25974 22513 26008 22529
rect 26042 22631 26108 22639
rect 26042 22597 26058 22631
rect 26092 22597 26108 22631
rect 26042 22563 26108 22597
rect 26042 22529 26058 22563
rect 26092 22529 26108 22563
rect 25874 22479 25890 22495
rect 25756 22461 25890 22479
rect 25924 22479 25940 22495
rect 26042 22495 26108 22529
rect 26142 22631 26202 22673
rect 26176 22597 26202 22631
rect 26142 22563 26202 22597
rect 26176 22529 26202 22563
rect 26142 22513 26202 22529
rect 26247 22593 26397 22637
rect 26247 22559 26259 22593
rect 26293 22559 26351 22593
rect 26385 22559 26397 22593
rect 26042 22479 26058 22495
rect 25924 22461 26058 22479
rect 26092 22479 26108 22495
rect 26247 22509 26397 22559
rect 26092 22466 26213 22479
rect 26092 22461 26158 22466
rect 25419 22445 26158 22461
rect 25419 22327 25488 22445
rect 25538 22402 26109 22411
rect 25538 22368 25546 22402
rect 26034 22395 26109 22402
rect 26034 22368 26058 22395
rect 25538 22361 25554 22368
rect 25588 22361 25638 22368
rect 25672 22361 25722 22368
rect 25756 22361 25806 22368
rect 25840 22361 25890 22368
rect 25924 22361 25974 22368
rect 26008 22361 26058 22368
rect 26092 22361 26109 22395
rect 26149 22327 26158 22445
rect 25419 22307 26158 22327
rect 25419 22289 25554 22307
rect 25538 22273 25554 22289
rect 25588 22289 25722 22307
rect 25588 22273 25604 22289
rect 25453 22239 25504 22255
rect 25453 22205 25470 22239
rect 25453 22163 25504 22205
rect 25538 22239 25604 22273
rect 25706 22273 25722 22289
rect 25756 22289 25890 22307
rect 25756 22273 25772 22289
rect 25538 22205 25554 22239
rect 25588 22205 25604 22239
rect 25538 22197 25604 22205
rect 25638 22239 25672 22255
rect 25638 22163 25672 22205
rect 25706 22239 25772 22273
rect 25874 22273 25890 22289
rect 25924 22289 26058 22307
rect 25924 22273 25940 22289
rect 25706 22205 25722 22239
rect 25756 22205 25772 22239
rect 25706 22197 25772 22205
rect 25806 22239 25840 22255
rect 25806 22163 25840 22205
rect 25874 22239 25940 22273
rect 26042 22273 26058 22289
rect 26092 22302 26158 22307
rect 26206 22302 26213 22466
rect 26247 22475 26259 22509
rect 26293 22475 26351 22509
rect 26385 22475 26397 22509
rect 26247 22440 26397 22475
rect 26092 22289 26213 22302
rect 26247 22291 26397 22308
rect 26092 22273 26108 22289
rect 25874 22205 25890 22239
rect 25924 22205 25940 22239
rect 25874 22197 25940 22205
rect 25974 22239 26008 22255
rect 25974 22163 26008 22205
rect 26042 22239 26108 22273
rect 26247 22257 26259 22291
rect 26293 22257 26351 22291
rect 26385 22257 26397 22291
rect 26042 22205 26058 22239
rect 26092 22205 26108 22239
rect 26042 22197 26108 22205
rect 26142 22239 26203 22255
rect 26176 22205 26203 22239
rect 26142 22163 26203 22205
rect 26247 22199 26397 22257
rect 25402 22129 25431 22163
rect 25465 22129 25523 22163
rect 25557 22129 25615 22163
rect 25649 22129 25707 22163
rect 25741 22129 25799 22163
rect 25833 22129 25891 22163
rect 25925 22129 25983 22163
rect 26017 22129 26075 22163
rect 26109 22129 26167 22163
rect 26201 22129 26259 22163
rect 26293 22129 26351 22163
rect 26385 22129 26414 22163
rect 24704 21928 24738 21990
rect 22340 21894 22436 21928
rect 24136 21898 24436 21928
rect 24136 21894 24232 21898
rect 24340 21894 24436 21898
rect 24642 21894 24738 21928
rect 12742 18819 13592 18832
rect 12742 18785 12871 18819
rect 13457 18785 13592 18819
rect 12742 18782 13592 18785
rect 12742 18722 12812 18782
rect 12742 18420 12775 18722
rect 12809 18420 12812 18722
rect 13512 18722 13592 18782
rect 12935 18682 12951 18716
rect 13119 18682 13135 18716
rect 13193 18682 13209 18716
rect 13377 18682 13393 18716
rect 12889 18632 12923 18639
rect 12742 18382 12812 18420
rect 12872 18623 12942 18632
rect 12872 18447 12889 18623
rect 12923 18462 12942 18623
rect 13147 18623 13181 18639
rect 13405 18632 13439 18639
rect 12923 18447 13072 18462
rect 12872 18382 13072 18447
rect 13392 18623 13452 18632
rect 13392 18462 13405 18623
rect 13147 18431 13181 18447
rect 13252 18447 13405 18462
rect 13439 18447 13452 18623
rect 13012 18302 13072 18382
rect 13252 18382 13452 18447
rect 13512 18420 13519 18722
rect 13553 18662 13592 18722
rect 25924 18689 26774 18702
rect 13553 18622 13792 18662
rect 13553 18442 13672 18622
rect 13772 18442 13792 18622
rect 13553 18420 13792 18442
rect 13512 18402 13792 18420
rect 25924 18655 26053 18689
rect 26639 18655 26774 18689
rect 25924 18652 26774 18655
rect 25924 18592 25994 18652
rect 13252 18302 13312 18382
rect 5716 18262 11260 18272
rect 5716 15582 5732 18262
rect 5772 18206 11212 18222
rect 5772 15632 5782 18206
rect 5980 17932 10996 17942
rect 5980 15912 5992 17932
rect 6032 17876 10942 17892
rect 6032 15962 6046 17876
rect 6906 17584 10642 17602
rect 6906 17514 6908 17584
rect 7340 17562 10642 17584
rect 10592 17522 10642 17562
rect 7340 17514 10642 17522
rect 6906 17482 10642 17514
rect 7506 17422 7540 17438
rect 7506 17230 7540 17246
rect 7764 17422 7798 17438
rect 7764 17230 7798 17246
rect 8022 17422 8056 17438
rect 8022 17230 8056 17246
rect 8280 17422 8314 17438
rect 8280 17230 8314 17246
rect 8538 17422 8572 17438
rect 8538 17230 8572 17246
rect 8796 17422 8830 17438
rect 8796 17230 8830 17246
rect 9054 17422 9088 17438
rect 9054 17230 9088 17246
rect 9312 17422 9346 17438
rect 9312 17230 9346 17246
rect 9570 17422 9604 17438
rect 9570 17230 9604 17246
rect 9828 17422 9862 17438
rect 9828 17230 9862 17246
rect 10086 17422 10120 17438
rect 10086 17230 10120 17246
rect 10344 17422 10378 17438
rect 10344 17230 10378 17246
rect 10602 17422 10636 17438
rect 10602 17230 10636 17246
rect 7552 17153 7568 17187
rect 7736 17153 7752 17187
rect 7810 17153 7826 17187
rect 7994 17153 8010 17187
rect 8068 17153 8084 17187
rect 8252 17153 8268 17187
rect 8326 17153 8342 17187
rect 8510 17153 8526 17187
rect 8584 17153 8600 17187
rect 8768 17153 8784 17187
rect 8842 17153 8858 17187
rect 9026 17153 9042 17187
rect 9100 17153 9116 17187
rect 9284 17153 9300 17187
rect 9358 17153 9374 17187
rect 9542 17153 9558 17187
rect 9616 17153 9632 17187
rect 9800 17153 9816 17187
rect 9874 17153 9890 17187
rect 10058 17153 10074 17187
rect 10132 17153 10148 17187
rect 10316 17153 10332 17187
rect 10390 17153 10406 17187
rect 10574 17153 10590 17187
rect 7810 17045 7826 17079
rect 7994 17045 8010 17079
rect 8584 17045 8600 17079
rect 8768 17045 8784 17079
rect 8842 17045 8858 17079
rect 9026 17045 9042 17079
rect 9616 17045 9632 17079
rect 9800 17045 9816 17079
rect 9874 17045 9890 17079
rect 10058 17045 10074 17079
rect 7506 16995 7540 17011
rect 7506 16803 7540 16819
rect 7764 16995 7798 17011
rect 7764 16803 7798 16819
rect 8022 16995 8056 17011
rect 8022 16803 8056 16819
rect 8280 16995 8314 17011
rect 8280 16803 8314 16819
rect 8538 16995 8572 17011
rect 8538 16803 8572 16819
rect 8796 16995 8830 17011
rect 8796 16803 8830 16819
rect 9054 16995 9088 17011
rect 9054 16803 9088 16819
rect 9312 16995 9346 17011
rect 9312 16803 9346 16819
rect 9570 16995 9604 17011
rect 9570 16803 9604 16819
rect 9828 16995 9862 17011
rect 9828 16803 9862 16819
rect 10086 16995 10120 17011
rect 10086 16803 10120 16819
rect 10344 16995 10378 17011
rect 10344 16803 10378 16819
rect 10602 16995 10636 17011
rect 10602 16803 10636 16819
rect 7552 16735 7568 16769
rect 7736 16735 7752 16769
rect 8068 16735 8084 16769
rect 8252 16735 8268 16769
rect 8326 16735 8342 16769
rect 8510 16735 8526 16769
rect 9100 16735 9116 16769
rect 9284 16735 9300 16769
rect 9358 16735 9374 16769
rect 9542 16735 9558 16769
rect 10132 16735 10148 16769
rect 10316 16735 10332 16769
rect 10390 16735 10406 16769
rect 10574 16735 10590 16769
rect 7552 16609 7568 16643
rect 7736 16609 7752 16643
rect 7810 16609 7826 16643
rect 7994 16609 8010 16643
rect 8068 16609 8084 16643
rect 8252 16609 8268 16643
rect 8326 16609 8342 16643
rect 8510 16609 8526 16643
rect 8584 16609 8600 16643
rect 8768 16609 8784 16643
rect 8842 16609 8858 16643
rect 9026 16609 9042 16643
rect 9100 16609 9116 16643
rect 9284 16609 9300 16643
rect 9358 16609 9374 16643
rect 9542 16609 9558 16643
rect 9616 16609 9632 16643
rect 9800 16609 9816 16643
rect 9874 16609 9890 16643
rect 10058 16609 10074 16643
rect 10132 16609 10148 16643
rect 10316 16609 10332 16643
rect 10390 16609 10406 16643
rect 10574 16609 10590 16643
rect 7506 16559 7540 16575
rect 7506 16483 7540 16499
rect 7764 16559 7798 16575
rect 7764 16483 7798 16499
rect 8022 16559 8056 16575
rect 8022 16483 8056 16499
rect 8280 16559 8314 16575
rect 8280 16483 8314 16499
rect 8538 16559 8572 16575
rect 8538 16483 8572 16499
rect 8796 16559 8830 16575
rect 8796 16483 8830 16499
rect 9054 16559 9088 16575
rect 9054 16483 9088 16499
rect 9312 16559 9346 16575
rect 9312 16483 9346 16499
rect 9570 16559 9604 16575
rect 9570 16483 9604 16499
rect 9828 16559 9862 16575
rect 9828 16483 9862 16499
rect 10086 16559 10120 16575
rect 10086 16483 10120 16499
rect 10344 16559 10378 16575
rect 10344 16483 10378 16499
rect 10602 16559 10636 16575
rect 10602 16483 10636 16499
rect 6906 16432 7392 16462
rect 6906 16422 6972 16432
rect 6906 16352 6908 16422
rect 6906 16342 6972 16352
rect 7372 16342 7392 16432
rect 6906 16322 7392 16342
rect 7502 16372 10642 16402
rect 7502 16322 7542 16372
rect 10592 16322 10642 16372
rect 7502 16292 10642 16322
rect 10930 15962 10942 17876
rect 6032 15952 10942 15962
rect 10982 15912 10996 17932
rect 5980 15896 10996 15912
rect 11194 15632 11212 18206
rect 5772 15622 11212 15632
rect 11252 15582 11260 18262
rect 13012 18222 13312 18302
rect 25924 18290 25957 18592
rect 25991 18290 25994 18592
rect 26694 18592 26774 18652
rect 26117 18552 26133 18586
rect 26301 18552 26317 18586
rect 26375 18552 26391 18586
rect 26559 18552 26575 18586
rect 26071 18502 26105 18509
rect 25924 18252 25994 18290
rect 26054 18493 26124 18502
rect 26054 18317 26071 18493
rect 26105 18332 26124 18493
rect 26329 18493 26363 18509
rect 26587 18502 26621 18509
rect 26105 18317 26254 18332
rect 26054 18252 26254 18317
rect 26574 18493 26634 18502
rect 26574 18332 26587 18493
rect 26329 18301 26363 18317
rect 26434 18317 26587 18332
rect 26621 18317 26634 18493
rect 12742 18155 12812 18182
rect 11508 18036 11604 18070
rect 11810 18036 11906 18070
rect 11508 17974 11542 18036
rect 11432 16382 11508 16402
rect 11872 17974 11906 18036
rect 11632 17940 11792 17942
rect 11632 17508 11638 17940
rect 11776 17508 11792 17940
rect 11632 17502 11792 17508
rect 11542 16382 11572 16402
rect 11432 15942 11452 16382
rect 11552 15942 11572 16382
rect 11432 15922 11508 15942
rect 5716 15566 11260 15582
rect 9532 15382 10692 15402
rect 9532 15376 9552 15382
rect 10672 15376 10692 15382
rect 9508 15302 9552 15376
rect 11304 15342 11400 15376
rect 10672 15302 10692 15342
rect 9508 15282 10692 15302
rect 11366 15302 11400 15342
rect 9508 15280 9542 15282
rect 11366 15280 11508 15302
rect 9508 15012 9542 15074
rect 11400 15074 11508 15280
rect 11542 15922 11572 15942
rect 11542 15074 11572 15302
rect 11366 15012 11572 15074
rect 12742 17861 12775 18155
rect 12809 17861 12812 18155
rect 12872 18127 12942 18182
rect 12872 17982 12889 18127
rect 12923 17982 12942 18127
rect 13112 18127 13212 18222
rect 12889 17935 12923 17951
rect 13112 17951 13147 18127
rect 13181 17951 13212 18127
rect 13392 18127 13452 18182
rect 13392 17982 13405 18127
rect 13112 17942 13212 17951
rect 13439 17982 13452 18127
rect 13512 18155 13792 18182
rect 13147 17935 13181 17942
rect 13405 17935 13439 17951
rect 12935 17867 12951 17901
rect 13119 17867 13135 17901
rect 13193 17867 13209 17901
rect 13377 17867 13393 17901
rect 12742 17802 12812 17861
rect 13512 17861 13519 18155
rect 13553 18142 13792 18155
rect 26194 18172 26254 18252
rect 26434 18252 26634 18317
rect 26694 18290 26701 18592
rect 26735 18532 26774 18592
rect 26735 18492 26974 18532
rect 26735 18312 26854 18492
rect 26954 18312 26974 18492
rect 26735 18290 26974 18312
rect 26694 18272 26974 18290
rect 26434 18172 26494 18252
rect 13553 17962 13672 18142
rect 13772 17962 13792 18142
rect 13553 17922 13792 17962
rect 18898 18132 24442 18142
rect 13553 17861 13592 17922
rect 13512 17802 13592 17861
rect 12742 17799 13592 17802
rect 12742 17765 12871 17799
rect 13457 17765 13592 17799
rect 12742 17732 13592 17765
rect 12742 17359 13592 17372
rect 12742 17325 12871 17359
rect 13457 17325 13592 17359
rect 12742 17322 13592 17325
rect 12742 17262 12812 17322
rect 12742 16960 12775 17262
rect 12809 16960 12812 17262
rect 13512 17262 13592 17322
rect 12935 17222 12951 17256
rect 13119 17222 13135 17256
rect 13193 17222 13209 17256
rect 13377 17222 13393 17256
rect 12889 17172 12923 17179
rect 12742 16922 12812 16960
rect 12872 17163 12942 17172
rect 12872 16987 12889 17163
rect 12923 17002 12942 17163
rect 13147 17163 13181 17179
rect 13405 17172 13439 17179
rect 12923 16987 13072 17002
rect 12872 16922 13072 16987
rect 13392 17163 13452 17172
rect 13392 17002 13405 17163
rect 13147 16971 13181 16987
rect 13252 16987 13405 17002
rect 13439 16987 13452 17163
rect 13012 16842 13072 16922
rect 13252 16922 13452 16987
rect 13512 16960 13519 17262
rect 13553 17202 13592 17262
rect 13553 17162 13792 17202
rect 13553 16982 13672 17162
rect 13772 16982 13792 17162
rect 13553 16960 13792 16982
rect 13512 16942 13792 16960
rect 13252 16842 13312 16922
rect 13012 16762 13312 16842
rect 12742 16695 12812 16722
rect 12742 16401 12775 16695
rect 12809 16401 12812 16695
rect 12872 16667 12942 16722
rect 12872 16522 12889 16667
rect 12923 16522 12942 16667
rect 13112 16667 13212 16762
rect 12889 16475 12923 16491
rect 13112 16491 13147 16667
rect 13181 16491 13212 16667
rect 13392 16667 13452 16722
rect 13392 16522 13405 16667
rect 13112 16482 13212 16491
rect 13439 16522 13452 16667
rect 13512 16695 13792 16722
rect 13147 16475 13181 16482
rect 13405 16475 13439 16491
rect 12935 16407 12951 16441
rect 13119 16407 13135 16441
rect 13193 16407 13209 16441
rect 13377 16407 13393 16441
rect 12742 16342 12812 16401
rect 13512 16401 13519 16695
rect 13553 16682 13792 16695
rect 13553 16502 13672 16682
rect 13772 16502 13792 16682
rect 13553 16462 13792 16502
rect 13553 16401 13592 16462
rect 13512 16342 13592 16401
rect 12742 16339 13592 16342
rect 12742 16305 12871 16339
rect 13457 16305 13592 16339
rect 12742 16272 13592 16305
rect 12570 15757 12599 15791
rect 12633 15757 12691 15791
rect 12725 15757 12783 15791
rect 12817 15757 12875 15791
rect 12909 15757 12967 15791
rect 13001 15757 13059 15791
rect 13093 15757 13151 15791
rect 13185 15757 13243 15791
rect 13277 15757 13335 15791
rect 13369 15757 13427 15791
rect 13461 15757 13519 15791
rect 13553 15757 13582 15791
rect 12621 15715 12672 15757
rect 12621 15681 12638 15715
rect 12621 15647 12672 15681
rect 12621 15613 12638 15647
rect 12621 15597 12672 15613
rect 12706 15715 12772 15723
rect 12706 15681 12722 15715
rect 12756 15681 12772 15715
rect 12706 15647 12772 15681
rect 12706 15613 12722 15647
rect 12756 15613 12772 15647
rect 12706 15579 12772 15613
rect 12806 15715 12840 15757
rect 12806 15647 12840 15681
rect 12806 15597 12840 15613
rect 12874 15715 12940 15723
rect 12874 15681 12890 15715
rect 12924 15681 12940 15715
rect 12874 15647 12940 15681
rect 12874 15613 12890 15647
rect 12924 15613 12940 15647
rect 12706 15563 12722 15579
rect 12587 15545 12722 15563
rect 12756 15563 12772 15579
rect 12874 15579 12940 15613
rect 12974 15715 13008 15757
rect 12974 15647 13008 15681
rect 12974 15597 13008 15613
rect 13042 15715 13108 15723
rect 13042 15681 13058 15715
rect 13092 15681 13108 15715
rect 13042 15647 13108 15681
rect 13042 15613 13058 15647
rect 13092 15613 13108 15647
rect 12874 15563 12890 15579
rect 12756 15545 12890 15563
rect 12924 15563 12940 15579
rect 13042 15579 13108 15613
rect 13142 15715 13176 15757
rect 13142 15647 13176 15681
rect 13142 15597 13176 15613
rect 13210 15715 13276 15723
rect 13210 15681 13226 15715
rect 13260 15681 13276 15715
rect 13210 15647 13276 15681
rect 13210 15613 13226 15647
rect 13260 15613 13276 15647
rect 13042 15563 13058 15579
rect 12924 15545 13058 15563
rect 13092 15563 13108 15579
rect 13210 15579 13276 15613
rect 13310 15715 13370 15757
rect 13344 15681 13370 15715
rect 13310 15647 13370 15681
rect 13344 15613 13370 15647
rect 13310 15597 13370 15613
rect 13415 15677 13565 15721
rect 13415 15643 13427 15677
rect 13461 15643 13519 15677
rect 13553 15643 13565 15677
rect 13210 15563 13226 15579
rect 13092 15545 13226 15563
rect 13260 15563 13276 15579
rect 13415 15593 13565 15643
rect 13260 15550 13381 15563
rect 13260 15545 13326 15550
rect 12587 15529 13326 15545
rect 12587 15411 12656 15529
rect 12706 15486 13277 15495
rect 12706 15452 12714 15486
rect 13202 15479 13277 15486
rect 13202 15452 13226 15479
rect 12706 15445 12722 15452
rect 12756 15445 12806 15452
rect 12840 15445 12890 15452
rect 12924 15445 12974 15452
rect 13008 15445 13058 15452
rect 13092 15445 13142 15452
rect 13176 15445 13226 15452
rect 13260 15445 13277 15479
rect 13317 15411 13326 15529
rect 12587 15391 13326 15411
rect 12587 15373 12722 15391
rect 12706 15357 12722 15373
rect 12756 15373 12890 15391
rect 12756 15357 12772 15373
rect 12621 15323 12672 15339
rect 12621 15289 12638 15323
rect 12621 15247 12672 15289
rect 12706 15323 12772 15357
rect 12874 15357 12890 15373
rect 12924 15373 13058 15391
rect 12924 15357 12940 15373
rect 12706 15289 12722 15323
rect 12756 15289 12772 15323
rect 12706 15281 12772 15289
rect 12806 15323 12840 15339
rect 12806 15247 12840 15289
rect 12874 15323 12940 15357
rect 13042 15357 13058 15373
rect 13092 15373 13226 15391
rect 13092 15357 13108 15373
rect 12874 15289 12890 15323
rect 12924 15289 12940 15323
rect 12874 15281 12940 15289
rect 12974 15323 13008 15339
rect 12974 15247 13008 15289
rect 13042 15323 13108 15357
rect 13210 15357 13226 15373
rect 13260 15386 13326 15391
rect 13374 15386 13381 15550
rect 13415 15559 13427 15593
rect 13461 15559 13519 15593
rect 13553 15559 13565 15593
rect 13415 15524 13565 15559
rect 18898 15452 18914 18132
rect 18954 18076 24394 18092
rect 18954 15502 18964 18076
rect 19162 17802 24178 17812
rect 19162 15782 19174 17802
rect 19214 17746 24124 17762
rect 19214 15832 19228 17746
rect 20088 17454 23824 17472
rect 20088 17384 20090 17454
rect 20522 17432 23824 17454
rect 23774 17392 23824 17432
rect 20522 17384 23824 17392
rect 20088 17352 23824 17384
rect 20688 17292 20722 17308
rect 20688 17100 20722 17116
rect 20946 17292 20980 17308
rect 20946 17100 20980 17116
rect 21204 17292 21238 17308
rect 21204 17100 21238 17116
rect 21462 17292 21496 17308
rect 21462 17100 21496 17116
rect 21720 17292 21754 17308
rect 21720 17100 21754 17116
rect 21978 17292 22012 17308
rect 21978 17100 22012 17116
rect 22236 17292 22270 17308
rect 22236 17100 22270 17116
rect 22494 17292 22528 17308
rect 22494 17100 22528 17116
rect 22752 17292 22786 17308
rect 22752 17100 22786 17116
rect 23010 17292 23044 17308
rect 23010 17100 23044 17116
rect 23268 17292 23302 17308
rect 23268 17100 23302 17116
rect 23526 17292 23560 17308
rect 23526 17100 23560 17116
rect 23784 17292 23818 17308
rect 23784 17100 23818 17116
rect 20734 17023 20750 17057
rect 20918 17023 20934 17057
rect 20992 17023 21008 17057
rect 21176 17023 21192 17057
rect 21250 17023 21266 17057
rect 21434 17023 21450 17057
rect 21508 17023 21524 17057
rect 21692 17023 21708 17057
rect 21766 17023 21782 17057
rect 21950 17023 21966 17057
rect 22024 17023 22040 17057
rect 22208 17023 22224 17057
rect 22282 17023 22298 17057
rect 22466 17023 22482 17057
rect 22540 17023 22556 17057
rect 22724 17023 22740 17057
rect 22798 17023 22814 17057
rect 22982 17023 22998 17057
rect 23056 17023 23072 17057
rect 23240 17023 23256 17057
rect 23314 17023 23330 17057
rect 23498 17023 23514 17057
rect 23572 17023 23588 17057
rect 23756 17023 23772 17057
rect 20992 16915 21008 16949
rect 21176 16915 21192 16949
rect 21766 16915 21782 16949
rect 21950 16915 21966 16949
rect 22024 16915 22040 16949
rect 22208 16915 22224 16949
rect 22798 16915 22814 16949
rect 22982 16915 22998 16949
rect 23056 16915 23072 16949
rect 23240 16915 23256 16949
rect 20688 16865 20722 16881
rect 20688 16673 20722 16689
rect 20946 16865 20980 16881
rect 20946 16673 20980 16689
rect 21204 16865 21238 16881
rect 21204 16673 21238 16689
rect 21462 16865 21496 16881
rect 21462 16673 21496 16689
rect 21720 16865 21754 16881
rect 21720 16673 21754 16689
rect 21978 16865 22012 16881
rect 21978 16673 22012 16689
rect 22236 16865 22270 16881
rect 22236 16673 22270 16689
rect 22494 16865 22528 16881
rect 22494 16673 22528 16689
rect 22752 16865 22786 16881
rect 22752 16673 22786 16689
rect 23010 16865 23044 16881
rect 23010 16673 23044 16689
rect 23268 16865 23302 16881
rect 23268 16673 23302 16689
rect 23526 16865 23560 16881
rect 23526 16673 23560 16689
rect 23784 16865 23818 16881
rect 23784 16673 23818 16689
rect 20734 16605 20750 16639
rect 20918 16605 20934 16639
rect 21250 16605 21266 16639
rect 21434 16605 21450 16639
rect 21508 16605 21524 16639
rect 21692 16605 21708 16639
rect 22282 16605 22298 16639
rect 22466 16605 22482 16639
rect 22540 16605 22556 16639
rect 22724 16605 22740 16639
rect 23314 16605 23330 16639
rect 23498 16605 23514 16639
rect 23572 16605 23588 16639
rect 23756 16605 23772 16639
rect 20734 16479 20750 16513
rect 20918 16479 20934 16513
rect 20992 16479 21008 16513
rect 21176 16479 21192 16513
rect 21250 16479 21266 16513
rect 21434 16479 21450 16513
rect 21508 16479 21524 16513
rect 21692 16479 21708 16513
rect 21766 16479 21782 16513
rect 21950 16479 21966 16513
rect 22024 16479 22040 16513
rect 22208 16479 22224 16513
rect 22282 16479 22298 16513
rect 22466 16479 22482 16513
rect 22540 16479 22556 16513
rect 22724 16479 22740 16513
rect 22798 16479 22814 16513
rect 22982 16479 22998 16513
rect 23056 16479 23072 16513
rect 23240 16479 23256 16513
rect 23314 16479 23330 16513
rect 23498 16479 23514 16513
rect 23572 16479 23588 16513
rect 23756 16479 23772 16513
rect 20688 16429 20722 16445
rect 20688 16353 20722 16369
rect 20946 16429 20980 16445
rect 20946 16353 20980 16369
rect 21204 16429 21238 16445
rect 21204 16353 21238 16369
rect 21462 16429 21496 16445
rect 21462 16353 21496 16369
rect 21720 16429 21754 16445
rect 21720 16353 21754 16369
rect 21978 16429 22012 16445
rect 21978 16353 22012 16369
rect 22236 16429 22270 16445
rect 22236 16353 22270 16369
rect 22494 16429 22528 16445
rect 22494 16353 22528 16369
rect 22752 16429 22786 16445
rect 22752 16353 22786 16369
rect 23010 16429 23044 16445
rect 23010 16353 23044 16369
rect 23268 16429 23302 16445
rect 23268 16353 23302 16369
rect 23526 16429 23560 16445
rect 23526 16353 23560 16369
rect 23784 16429 23818 16445
rect 23784 16353 23818 16369
rect 20088 16302 20574 16332
rect 20088 16292 20154 16302
rect 20088 16222 20090 16292
rect 20088 16212 20154 16222
rect 20554 16212 20574 16302
rect 20088 16192 20574 16212
rect 20684 16242 23824 16272
rect 20684 16192 20724 16242
rect 23774 16192 23824 16242
rect 20684 16162 23824 16192
rect 24112 15832 24124 17746
rect 19214 15822 24124 15832
rect 24164 15782 24178 17802
rect 19162 15766 24178 15782
rect 24376 15502 24394 18076
rect 18954 15492 24394 15502
rect 24434 15452 24442 18132
rect 26194 18092 26494 18172
rect 25924 18025 25994 18052
rect 24690 17906 24786 17940
rect 24992 17906 25088 17940
rect 24690 17844 24724 17906
rect 24614 16252 24690 16272
rect 25054 17844 25088 17906
rect 24814 17810 24974 17812
rect 24814 17378 24820 17810
rect 24958 17378 24974 17810
rect 24814 17372 24974 17378
rect 24724 16252 24754 16272
rect 24614 15812 24634 16252
rect 24734 15812 24754 16252
rect 24614 15792 24690 15812
rect 18898 15436 24442 15452
rect 13260 15373 13381 15386
rect 13415 15375 13565 15392
rect 13260 15357 13276 15373
rect 13042 15289 13058 15323
rect 13092 15289 13108 15323
rect 13042 15281 13108 15289
rect 13142 15323 13176 15339
rect 13142 15247 13176 15289
rect 13210 15323 13276 15357
rect 13415 15341 13427 15375
rect 13461 15341 13519 15375
rect 13553 15341 13565 15375
rect 13210 15289 13226 15323
rect 13260 15289 13276 15323
rect 13210 15281 13276 15289
rect 13310 15323 13371 15339
rect 13344 15289 13371 15323
rect 13310 15247 13371 15289
rect 13415 15283 13565 15341
rect 22714 15252 23874 15272
rect 12570 15213 12599 15247
rect 12633 15213 12691 15247
rect 12725 15213 12783 15247
rect 12817 15213 12875 15247
rect 12909 15213 12967 15247
rect 13001 15213 13059 15247
rect 13093 15213 13151 15247
rect 13185 15213 13243 15247
rect 13277 15213 13335 15247
rect 13369 15213 13427 15247
rect 13461 15213 13519 15247
rect 13553 15213 13582 15247
rect 22714 15246 22734 15252
rect 23854 15246 23874 15252
rect 11872 15012 11906 15074
rect 9508 14978 9604 15012
rect 11304 14982 11604 15012
rect 11304 14978 11400 14982
rect 11508 14978 11604 14982
rect 11810 14978 11906 15012
rect 22690 15172 22734 15246
rect 24486 15212 24582 15246
rect 23854 15172 23874 15212
rect 22690 15152 23874 15172
rect 24548 15172 24582 15212
rect 22690 15150 22724 15152
rect 24548 15150 24690 15172
rect 22690 14882 22724 14944
rect 24582 14944 24690 15150
rect 24724 15792 24754 15812
rect 24724 14944 24754 15172
rect 24548 14882 24754 14944
rect 25924 17731 25957 18025
rect 25991 17731 25994 18025
rect 26054 17997 26124 18052
rect 26054 17852 26071 17997
rect 26105 17852 26124 17997
rect 26294 17997 26394 18092
rect 26071 17805 26105 17821
rect 26294 17821 26329 17997
rect 26363 17821 26394 17997
rect 26574 17997 26634 18052
rect 26574 17852 26587 17997
rect 26294 17812 26394 17821
rect 26621 17852 26634 17997
rect 26694 18025 26974 18052
rect 26329 17805 26363 17812
rect 26587 17805 26621 17821
rect 26117 17737 26133 17771
rect 26301 17737 26317 17771
rect 26375 17737 26391 17771
rect 26559 17737 26575 17771
rect 25924 17672 25994 17731
rect 26694 17731 26701 18025
rect 26735 18012 26974 18025
rect 26735 17832 26854 18012
rect 26954 17832 26974 18012
rect 26735 17792 26974 17832
rect 26735 17731 26774 17792
rect 26694 17672 26774 17731
rect 25924 17669 26774 17672
rect 25924 17635 26053 17669
rect 26639 17635 26774 17669
rect 25924 17602 26774 17635
rect 25924 17229 26774 17242
rect 25924 17195 26053 17229
rect 26639 17195 26774 17229
rect 25924 17192 26774 17195
rect 25924 17132 25994 17192
rect 25924 16830 25957 17132
rect 25991 16830 25994 17132
rect 26694 17132 26774 17192
rect 26117 17092 26133 17126
rect 26301 17092 26317 17126
rect 26375 17092 26391 17126
rect 26559 17092 26575 17126
rect 26071 17042 26105 17049
rect 25924 16792 25994 16830
rect 26054 17033 26124 17042
rect 26054 16857 26071 17033
rect 26105 16872 26124 17033
rect 26329 17033 26363 17049
rect 26587 17042 26621 17049
rect 26105 16857 26254 16872
rect 26054 16792 26254 16857
rect 26574 17033 26634 17042
rect 26574 16872 26587 17033
rect 26329 16841 26363 16857
rect 26434 16857 26587 16872
rect 26621 16857 26634 17033
rect 26194 16712 26254 16792
rect 26434 16792 26634 16857
rect 26694 16830 26701 17132
rect 26735 17072 26774 17132
rect 26735 17032 26974 17072
rect 26735 16852 26854 17032
rect 26954 16852 26974 17032
rect 26735 16830 26974 16852
rect 26694 16812 26974 16830
rect 26434 16712 26494 16792
rect 26194 16632 26494 16712
rect 25924 16565 25994 16592
rect 25924 16271 25957 16565
rect 25991 16271 25994 16565
rect 26054 16537 26124 16592
rect 26054 16392 26071 16537
rect 26105 16392 26124 16537
rect 26294 16537 26394 16632
rect 26071 16345 26105 16361
rect 26294 16361 26329 16537
rect 26363 16361 26394 16537
rect 26574 16537 26634 16592
rect 26574 16392 26587 16537
rect 26294 16352 26394 16361
rect 26621 16392 26634 16537
rect 26694 16565 26974 16592
rect 26329 16345 26363 16352
rect 26587 16345 26621 16361
rect 26117 16277 26133 16311
rect 26301 16277 26317 16311
rect 26375 16277 26391 16311
rect 26559 16277 26575 16311
rect 25924 16212 25994 16271
rect 26694 16271 26701 16565
rect 26735 16552 26974 16565
rect 26735 16372 26854 16552
rect 26954 16372 26974 16552
rect 26735 16332 26974 16372
rect 26735 16271 26774 16332
rect 26694 16212 26774 16271
rect 25924 16209 26774 16212
rect 25924 16175 26053 16209
rect 26639 16175 26774 16209
rect 25924 16142 26774 16175
rect 25752 15627 25781 15661
rect 25815 15627 25873 15661
rect 25907 15627 25965 15661
rect 25999 15627 26057 15661
rect 26091 15627 26149 15661
rect 26183 15627 26241 15661
rect 26275 15627 26333 15661
rect 26367 15627 26425 15661
rect 26459 15627 26517 15661
rect 26551 15627 26609 15661
rect 26643 15627 26701 15661
rect 26735 15627 26764 15661
rect 25803 15585 25854 15627
rect 25803 15551 25820 15585
rect 25803 15517 25854 15551
rect 25803 15483 25820 15517
rect 25803 15467 25854 15483
rect 25888 15585 25954 15593
rect 25888 15551 25904 15585
rect 25938 15551 25954 15585
rect 25888 15517 25954 15551
rect 25888 15483 25904 15517
rect 25938 15483 25954 15517
rect 25888 15449 25954 15483
rect 25988 15585 26022 15627
rect 25988 15517 26022 15551
rect 25988 15467 26022 15483
rect 26056 15585 26122 15593
rect 26056 15551 26072 15585
rect 26106 15551 26122 15585
rect 26056 15517 26122 15551
rect 26056 15483 26072 15517
rect 26106 15483 26122 15517
rect 25888 15433 25904 15449
rect 25769 15415 25904 15433
rect 25938 15433 25954 15449
rect 26056 15449 26122 15483
rect 26156 15585 26190 15627
rect 26156 15517 26190 15551
rect 26156 15467 26190 15483
rect 26224 15585 26290 15593
rect 26224 15551 26240 15585
rect 26274 15551 26290 15585
rect 26224 15517 26290 15551
rect 26224 15483 26240 15517
rect 26274 15483 26290 15517
rect 26056 15433 26072 15449
rect 25938 15415 26072 15433
rect 26106 15433 26122 15449
rect 26224 15449 26290 15483
rect 26324 15585 26358 15627
rect 26324 15517 26358 15551
rect 26324 15467 26358 15483
rect 26392 15585 26458 15593
rect 26392 15551 26408 15585
rect 26442 15551 26458 15585
rect 26392 15517 26458 15551
rect 26392 15483 26408 15517
rect 26442 15483 26458 15517
rect 26224 15433 26240 15449
rect 26106 15415 26240 15433
rect 26274 15433 26290 15449
rect 26392 15449 26458 15483
rect 26492 15585 26552 15627
rect 26526 15551 26552 15585
rect 26492 15517 26552 15551
rect 26526 15483 26552 15517
rect 26492 15467 26552 15483
rect 26597 15547 26747 15591
rect 26597 15513 26609 15547
rect 26643 15513 26701 15547
rect 26735 15513 26747 15547
rect 26392 15433 26408 15449
rect 26274 15415 26408 15433
rect 26442 15433 26458 15449
rect 26597 15463 26747 15513
rect 26442 15420 26563 15433
rect 26442 15415 26508 15420
rect 25769 15399 26508 15415
rect 25769 15281 25838 15399
rect 25888 15356 26459 15365
rect 25888 15322 25896 15356
rect 26384 15349 26459 15356
rect 26384 15322 26408 15349
rect 25888 15315 25904 15322
rect 25938 15315 25988 15322
rect 26022 15315 26072 15322
rect 26106 15315 26156 15322
rect 26190 15315 26240 15322
rect 26274 15315 26324 15322
rect 26358 15315 26408 15322
rect 26442 15315 26459 15349
rect 26499 15281 26508 15399
rect 25769 15261 26508 15281
rect 25769 15243 25904 15261
rect 25888 15227 25904 15243
rect 25938 15243 26072 15261
rect 25938 15227 25954 15243
rect 25803 15193 25854 15209
rect 25803 15159 25820 15193
rect 25803 15117 25854 15159
rect 25888 15193 25954 15227
rect 26056 15227 26072 15243
rect 26106 15243 26240 15261
rect 26106 15227 26122 15243
rect 25888 15159 25904 15193
rect 25938 15159 25954 15193
rect 25888 15151 25954 15159
rect 25988 15193 26022 15209
rect 25988 15117 26022 15159
rect 26056 15193 26122 15227
rect 26224 15227 26240 15243
rect 26274 15243 26408 15261
rect 26274 15227 26290 15243
rect 26056 15159 26072 15193
rect 26106 15159 26122 15193
rect 26056 15151 26122 15159
rect 26156 15193 26190 15209
rect 26156 15117 26190 15159
rect 26224 15193 26290 15227
rect 26392 15227 26408 15243
rect 26442 15256 26508 15261
rect 26556 15256 26563 15420
rect 26597 15429 26609 15463
rect 26643 15429 26701 15463
rect 26735 15429 26747 15463
rect 26597 15394 26747 15429
rect 26442 15243 26563 15256
rect 26597 15245 26747 15262
rect 26442 15227 26458 15243
rect 26224 15159 26240 15193
rect 26274 15159 26290 15193
rect 26224 15151 26290 15159
rect 26324 15193 26358 15209
rect 26324 15117 26358 15159
rect 26392 15193 26458 15227
rect 26597 15211 26609 15245
rect 26643 15211 26701 15245
rect 26735 15211 26747 15245
rect 26392 15159 26408 15193
rect 26442 15159 26458 15193
rect 26392 15151 26458 15159
rect 26492 15193 26553 15209
rect 26526 15159 26553 15193
rect 26492 15117 26553 15159
rect 26597 15153 26747 15211
rect 25752 15083 25781 15117
rect 25815 15083 25873 15117
rect 25907 15083 25965 15117
rect 25999 15083 26057 15117
rect 26091 15083 26149 15117
rect 26183 15083 26241 15117
rect 26275 15083 26333 15117
rect 26367 15083 26425 15117
rect 26459 15083 26517 15117
rect 26551 15083 26609 15117
rect 26643 15083 26701 15117
rect 26735 15083 26764 15117
rect 25054 14882 25088 14944
rect 22690 14848 22786 14882
rect 24486 14852 24786 14882
rect 24486 14848 24582 14852
rect 24690 14848 24786 14852
rect 24992 14848 25088 14882
<< viali >>
rect 12935 38358 13103 38392
rect 13193 38358 13361 38392
rect 12873 38123 12907 38299
rect 13131 38123 13165 38299
rect 13389 38123 13423 38299
rect 13656 38118 13756 38298
rect 25723 38476 25891 38510
rect 25981 38476 26149 38510
rect 25661 38241 25695 38417
rect 25919 38241 25953 38417
rect 26177 38241 26211 38417
rect 26444 38236 26544 38416
rect 5716 37898 5766 37938
rect 5766 37898 11166 37938
rect 11166 37898 11236 37938
rect 5716 37858 5756 37898
rect 5716 35328 5756 37858
rect 5716 35298 5756 35328
rect 5976 37568 6036 37608
rect 6036 37568 10886 37608
rect 10886 37568 10966 37608
rect 5976 37538 6016 37568
rect 5976 35668 6016 37538
rect 5976 35628 6016 35668
rect 6996 37198 7324 37238
rect 7324 37198 7566 37238
rect 7566 37198 10576 37238
rect 7490 36922 7524 37098
rect 7748 36922 7782 37098
rect 8006 36922 8040 37098
rect 8264 36922 8298 37098
rect 8522 36922 8556 37098
rect 8780 36922 8814 37098
rect 9038 36922 9072 37098
rect 9296 36922 9330 37098
rect 9554 36922 9588 37098
rect 9812 36922 9846 37098
rect 10070 36922 10104 37098
rect 10328 36922 10362 37098
rect 10586 36922 10620 37098
rect 7552 36829 7720 36863
rect 7810 36829 7978 36863
rect 8068 36829 8236 36863
rect 8326 36829 8494 36863
rect 8584 36829 8752 36863
rect 8842 36829 9010 36863
rect 9100 36829 9268 36863
rect 9358 36829 9526 36863
rect 9616 36829 9784 36863
rect 9874 36829 10042 36863
rect 10132 36829 10300 36863
rect 10390 36829 10558 36863
rect 7810 36721 7978 36755
rect 8584 36721 8752 36755
rect 8842 36721 9010 36755
rect 9616 36721 9784 36755
rect 9874 36721 10042 36755
rect 7490 36495 7524 36671
rect 7748 36495 7782 36671
rect 8006 36495 8040 36671
rect 8264 36495 8298 36671
rect 8522 36495 8556 36671
rect 8780 36495 8814 36671
rect 9038 36495 9072 36671
rect 9296 36495 9330 36671
rect 9554 36495 9588 36671
rect 9812 36495 9846 36671
rect 10070 36495 10104 36671
rect 10328 36495 10362 36671
rect 10586 36495 10620 36671
rect 7552 36411 7720 36445
rect 8068 36411 8236 36445
rect 8326 36411 8494 36445
rect 9100 36411 9268 36445
rect 9358 36411 9526 36445
rect 10132 36411 10300 36445
rect 10390 36411 10558 36445
rect 7552 36285 7720 36319
rect 7810 36285 7978 36319
rect 8068 36285 8236 36319
rect 8326 36285 8494 36319
rect 8584 36285 8752 36319
rect 8842 36285 9010 36319
rect 9100 36285 9268 36319
rect 9358 36285 9526 36319
rect 9616 36285 9784 36319
rect 9874 36285 10042 36319
rect 10132 36285 10300 36319
rect 10390 36285 10558 36319
rect 7490 36175 7524 36235
rect 7748 36175 7782 36235
rect 8006 36175 8040 36235
rect 8264 36175 8298 36235
rect 8522 36175 8556 36235
rect 8780 36175 8814 36235
rect 9038 36175 9072 36235
rect 9296 36175 9330 36235
rect 9554 36175 9588 36235
rect 9812 36175 9846 36235
rect 10070 36175 10104 36235
rect 10328 36175 10362 36235
rect 10586 36175 10620 36235
rect 6956 36098 7356 36108
rect 6956 36028 7324 36098
rect 7324 36028 7356 36098
rect 6956 36018 7356 36028
rect 7526 35998 10576 36048
rect 10926 37548 10966 37568
rect 10926 35658 10966 37548
rect 10926 35628 10966 35658
rect 5976 35588 6036 35628
rect 6036 35588 10896 35628
rect 10896 35588 10966 35628
rect 11196 37868 11236 37898
rect 11196 35318 11236 37868
rect 11196 35298 11236 35318
rect 5716 35258 5796 35298
rect 5796 35258 11166 35298
rect 11166 35258 11236 35298
rect 11636 37198 11756 37598
rect 12873 37627 12907 37803
rect 13131 37627 13165 37803
rect 13389 37627 13423 37803
rect 12935 37543 13103 37577
rect 13193 37543 13361 37577
rect 13656 37638 13756 37818
rect 12935 36898 13103 36932
rect 13193 36898 13361 36932
rect 12873 36663 12907 36839
rect 13131 36663 13165 36839
rect 13389 36663 13423 36839
rect 13656 36658 13756 36838
rect 12873 36167 12907 36343
rect 13131 36167 13165 36343
rect 13389 36167 13423 36343
rect 12935 36083 13103 36117
rect 13193 36083 13361 36117
rect 13656 36178 13756 36358
rect 12583 35433 12617 35467
rect 12675 35433 12709 35467
rect 12767 35433 12801 35467
rect 12859 35433 12893 35467
rect 12951 35433 12985 35467
rect 13043 35433 13077 35467
rect 13135 35433 13169 35467
rect 13227 35433 13261 35467
rect 13319 35433 13353 35467
rect 13411 35433 13445 35467
rect 13503 35433 13537 35467
rect 18504 38016 18554 38056
rect 18554 38016 23954 38056
rect 23954 38016 24024 38056
rect 18504 37976 18544 38016
rect 18504 35446 18544 37976
rect 18504 35416 18544 35446
rect 18764 37686 18824 37726
rect 18824 37686 23674 37726
rect 23674 37686 23754 37726
rect 18764 37656 18804 37686
rect 18764 35786 18804 37656
rect 18764 35746 18804 35786
rect 19784 37316 20112 37356
rect 20112 37316 20354 37356
rect 20354 37316 23364 37356
rect 20278 37040 20312 37216
rect 20536 37040 20570 37216
rect 20794 37040 20828 37216
rect 21052 37040 21086 37216
rect 21310 37040 21344 37216
rect 21568 37040 21602 37216
rect 21826 37040 21860 37216
rect 22084 37040 22118 37216
rect 22342 37040 22376 37216
rect 22600 37040 22634 37216
rect 22858 37040 22892 37216
rect 23116 37040 23150 37216
rect 23374 37040 23408 37216
rect 20340 36947 20508 36981
rect 20598 36947 20766 36981
rect 20856 36947 21024 36981
rect 21114 36947 21282 36981
rect 21372 36947 21540 36981
rect 21630 36947 21798 36981
rect 21888 36947 22056 36981
rect 22146 36947 22314 36981
rect 22404 36947 22572 36981
rect 22662 36947 22830 36981
rect 22920 36947 23088 36981
rect 23178 36947 23346 36981
rect 20598 36839 20766 36873
rect 21372 36839 21540 36873
rect 21630 36839 21798 36873
rect 22404 36839 22572 36873
rect 22662 36839 22830 36873
rect 20278 36613 20312 36789
rect 20536 36613 20570 36789
rect 20794 36613 20828 36789
rect 21052 36613 21086 36789
rect 21310 36613 21344 36789
rect 21568 36613 21602 36789
rect 21826 36613 21860 36789
rect 22084 36613 22118 36789
rect 22342 36613 22376 36789
rect 22600 36613 22634 36789
rect 22858 36613 22892 36789
rect 23116 36613 23150 36789
rect 23374 36613 23408 36789
rect 20340 36529 20508 36563
rect 20856 36529 21024 36563
rect 21114 36529 21282 36563
rect 21888 36529 22056 36563
rect 22146 36529 22314 36563
rect 22920 36529 23088 36563
rect 23178 36529 23346 36563
rect 20340 36403 20508 36437
rect 20598 36403 20766 36437
rect 20856 36403 21024 36437
rect 21114 36403 21282 36437
rect 21372 36403 21540 36437
rect 21630 36403 21798 36437
rect 21888 36403 22056 36437
rect 22146 36403 22314 36437
rect 22404 36403 22572 36437
rect 22662 36403 22830 36437
rect 22920 36403 23088 36437
rect 23178 36403 23346 36437
rect 20278 36293 20312 36353
rect 20536 36293 20570 36353
rect 20794 36293 20828 36353
rect 21052 36293 21086 36353
rect 21310 36293 21344 36353
rect 21568 36293 21602 36353
rect 21826 36293 21860 36353
rect 22084 36293 22118 36353
rect 22342 36293 22376 36353
rect 22600 36293 22634 36353
rect 22858 36293 22892 36353
rect 23116 36293 23150 36353
rect 23374 36293 23408 36353
rect 19744 36216 20144 36226
rect 19744 36146 20112 36216
rect 20112 36146 20144 36216
rect 19744 36136 20144 36146
rect 20314 36116 23364 36166
rect 23714 37666 23754 37686
rect 23714 35776 23754 37666
rect 23714 35746 23754 35776
rect 18764 35706 18824 35746
rect 18824 35706 23684 35746
rect 23684 35706 23754 35746
rect 23984 37986 24024 38016
rect 23984 35436 24024 37986
rect 23984 35416 24024 35436
rect 18504 35376 18584 35416
rect 18584 35376 23954 35416
rect 23954 35376 24024 35416
rect 24424 37316 24544 37716
rect 24224 35736 24280 36176
rect 24280 35736 24314 36176
rect 24314 35736 24324 36176
rect 12698 35155 13186 35162
rect 12698 35128 12706 35155
rect 12706 35128 12740 35155
rect 12740 35128 12790 35155
rect 12790 35128 12824 35155
rect 12824 35128 12874 35155
rect 12874 35128 12908 35155
rect 12908 35128 12958 35155
rect 12958 35128 12992 35155
rect 12992 35128 13042 35155
rect 13042 35128 13076 35155
rect 13076 35128 13126 35155
rect 13126 35128 13160 35155
rect 13160 35128 13186 35155
rect 13310 35062 13358 35226
rect 22324 35170 23444 35176
rect 22324 35136 22376 35170
rect 22376 35136 23444 35170
rect 22324 35096 23444 35136
rect 12583 34889 12617 34923
rect 12675 34889 12709 34923
rect 12767 34889 12801 34923
rect 12859 34889 12893 34923
rect 12951 34889 12985 34923
rect 13043 34889 13077 34923
rect 13135 34889 13169 34923
rect 13227 34889 13261 34923
rect 13319 34889 13353 34923
rect 13411 34889 13445 34923
rect 13503 34889 13537 34923
rect 22428 34918 22825 35024
rect 23627 34918 24024 35024
rect 24426 34920 24532 35317
rect 25661 37745 25695 37921
rect 25919 37745 25953 37921
rect 26177 37745 26211 37921
rect 25723 37661 25891 37695
rect 25981 37661 26149 37695
rect 26444 37756 26544 37936
rect 25723 37016 25891 37050
rect 25981 37016 26149 37050
rect 25661 36781 25695 36957
rect 25919 36781 25953 36957
rect 26177 36781 26211 36957
rect 26444 36776 26544 36956
rect 25661 36285 25695 36461
rect 25919 36285 25953 36461
rect 26177 36285 26211 36461
rect 25723 36201 25891 36235
rect 25981 36201 26149 36235
rect 26444 36296 26544 36476
rect 25371 35551 25405 35585
rect 25463 35551 25497 35585
rect 25555 35551 25589 35585
rect 25647 35551 25681 35585
rect 25739 35551 25773 35585
rect 25831 35551 25865 35585
rect 25923 35551 25957 35585
rect 26015 35551 26049 35585
rect 26107 35551 26141 35585
rect 26199 35551 26233 35585
rect 26291 35551 26325 35585
rect 25486 35273 25974 35280
rect 25486 35246 25494 35273
rect 25494 35246 25528 35273
rect 25528 35246 25578 35273
rect 25578 35246 25612 35273
rect 25612 35246 25662 35273
rect 25662 35246 25696 35273
rect 25696 35246 25746 35273
rect 25746 35246 25780 35273
rect 25780 35246 25830 35273
rect 25830 35246 25864 35273
rect 25864 35246 25914 35273
rect 25914 35246 25948 35273
rect 25948 35246 25974 35273
rect 26098 35180 26146 35344
rect 25371 35007 25405 35041
rect 25463 35007 25497 35041
rect 25555 35007 25589 35041
rect 25647 35007 25681 35041
rect 25739 35007 25773 35041
rect 25831 35007 25865 35041
rect 25923 35007 25957 35041
rect 26015 35007 26049 35041
rect 26107 35007 26141 35041
rect 26199 35007 26233 35041
rect 26291 35007 26325 35041
rect 12955 32432 13123 32466
rect 13213 32432 13381 32466
rect 12893 32197 12927 32373
rect 13151 32197 13185 32373
rect 13409 32197 13443 32373
rect 13676 32192 13776 32372
rect 25687 32356 25855 32390
rect 25945 32356 26113 32390
rect 25625 32121 25659 32297
rect 25883 32121 25917 32297
rect 26141 32121 26175 32297
rect 5736 31972 5786 32012
rect 5786 31972 11186 32012
rect 11186 31972 11256 32012
rect 5736 31932 5776 31972
rect 5736 29402 5776 31932
rect 5736 29372 5776 29402
rect 5996 31642 6056 31682
rect 6056 31642 10906 31682
rect 10906 31642 10986 31682
rect 5996 31612 6036 31642
rect 5996 29742 6036 31612
rect 5996 29702 6036 29742
rect 7016 31272 7344 31312
rect 7344 31272 7586 31312
rect 7586 31272 10596 31312
rect 7510 30996 7544 31172
rect 7768 30996 7802 31172
rect 8026 30996 8060 31172
rect 8284 30996 8318 31172
rect 8542 30996 8576 31172
rect 8800 30996 8834 31172
rect 9058 30996 9092 31172
rect 9316 30996 9350 31172
rect 9574 30996 9608 31172
rect 9832 30996 9866 31172
rect 10090 30996 10124 31172
rect 10348 30996 10382 31172
rect 10606 30996 10640 31172
rect 7572 30903 7740 30937
rect 7830 30903 7998 30937
rect 8088 30903 8256 30937
rect 8346 30903 8514 30937
rect 8604 30903 8772 30937
rect 8862 30903 9030 30937
rect 9120 30903 9288 30937
rect 9378 30903 9546 30937
rect 9636 30903 9804 30937
rect 9894 30903 10062 30937
rect 10152 30903 10320 30937
rect 10410 30903 10578 30937
rect 7830 30795 7998 30829
rect 8604 30795 8772 30829
rect 8862 30795 9030 30829
rect 9636 30795 9804 30829
rect 9894 30795 10062 30829
rect 7510 30569 7544 30745
rect 7768 30569 7802 30745
rect 8026 30569 8060 30745
rect 8284 30569 8318 30745
rect 8542 30569 8576 30745
rect 8800 30569 8834 30745
rect 9058 30569 9092 30745
rect 9316 30569 9350 30745
rect 9574 30569 9608 30745
rect 9832 30569 9866 30745
rect 10090 30569 10124 30745
rect 10348 30569 10382 30745
rect 10606 30569 10640 30745
rect 7572 30485 7740 30519
rect 8088 30485 8256 30519
rect 8346 30485 8514 30519
rect 9120 30485 9288 30519
rect 9378 30485 9546 30519
rect 10152 30485 10320 30519
rect 10410 30485 10578 30519
rect 7572 30359 7740 30393
rect 7830 30359 7998 30393
rect 8088 30359 8256 30393
rect 8346 30359 8514 30393
rect 8604 30359 8772 30393
rect 8862 30359 9030 30393
rect 9120 30359 9288 30393
rect 9378 30359 9546 30393
rect 9636 30359 9804 30393
rect 9894 30359 10062 30393
rect 10152 30359 10320 30393
rect 10410 30359 10578 30393
rect 7510 30249 7544 30309
rect 7768 30249 7802 30309
rect 8026 30249 8060 30309
rect 8284 30249 8318 30309
rect 8542 30249 8576 30309
rect 8800 30249 8834 30309
rect 9058 30249 9092 30309
rect 9316 30249 9350 30309
rect 9574 30249 9608 30309
rect 9832 30249 9866 30309
rect 10090 30249 10124 30309
rect 10348 30249 10382 30309
rect 10606 30249 10640 30309
rect 6976 30172 7376 30182
rect 6976 30102 7344 30172
rect 7344 30102 7376 30172
rect 6976 30092 7376 30102
rect 7546 30072 10596 30122
rect 10946 31622 10986 31642
rect 10946 29732 10986 31622
rect 10946 29702 10986 29732
rect 5996 29662 6056 29702
rect 6056 29662 10916 29702
rect 10916 29662 10986 29702
rect 11216 31942 11256 31972
rect 11216 29392 11256 31942
rect 11216 29372 11256 29392
rect 5736 29332 5816 29372
rect 5816 29332 11186 29372
rect 11186 29332 11256 29372
rect 26408 32116 26508 32296
rect 11656 31272 11776 31672
rect 11456 29692 11512 30132
rect 11512 29692 11546 30132
rect 11546 29692 11556 30132
rect 9556 29126 10676 29132
rect 9556 29092 9608 29126
rect 9608 29092 10676 29126
rect 9556 29052 10676 29092
rect 9660 28874 10057 28980
rect 10859 28874 11256 28980
rect 11658 28876 11764 29273
rect 12893 31701 12927 31877
rect 13151 31701 13185 31877
rect 13409 31701 13443 31877
rect 12955 31617 13123 31651
rect 13213 31617 13381 31651
rect 13676 31712 13776 31892
rect 12955 30972 13123 31006
rect 13213 30972 13381 31006
rect 12893 30737 12927 30913
rect 13151 30737 13185 30913
rect 13409 30737 13443 30913
rect 13676 30732 13776 30912
rect 12893 30241 12927 30417
rect 13151 30241 13185 30417
rect 13409 30241 13443 30417
rect 12955 30157 13123 30191
rect 13213 30157 13381 30191
rect 13676 30252 13776 30432
rect 12603 29507 12637 29541
rect 12695 29507 12729 29541
rect 12787 29507 12821 29541
rect 12879 29507 12913 29541
rect 12971 29507 13005 29541
rect 13063 29507 13097 29541
rect 13155 29507 13189 29541
rect 13247 29507 13281 29541
rect 13339 29507 13373 29541
rect 13431 29507 13465 29541
rect 13523 29507 13557 29541
rect 12718 29229 13206 29236
rect 12718 29202 12726 29229
rect 12726 29202 12760 29229
rect 12760 29202 12810 29229
rect 12810 29202 12844 29229
rect 12844 29202 12894 29229
rect 12894 29202 12928 29229
rect 12928 29202 12978 29229
rect 12978 29202 13012 29229
rect 13012 29202 13062 29229
rect 13062 29202 13096 29229
rect 13096 29202 13146 29229
rect 13146 29202 13180 29229
rect 13180 29202 13206 29229
rect 13330 29136 13378 29300
rect 18468 31896 18518 31936
rect 18518 31896 23918 31936
rect 23918 31896 23988 31936
rect 18468 31856 18508 31896
rect 18468 29326 18508 31856
rect 18468 29296 18508 29326
rect 18728 31566 18788 31606
rect 18788 31566 23638 31606
rect 23638 31566 23718 31606
rect 18728 31536 18768 31566
rect 18728 29666 18768 31536
rect 18728 29626 18768 29666
rect 19748 31196 20076 31236
rect 20076 31196 20318 31236
rect 20318 31196 23328 31236
rect 20242 30920 20276 31096
rect 20500 30920 20534 31096
rect 20758 30920 20792 31096
rect 21016 30920 21050 31096
rect 21274 30920 21308 31096
rect 21532 30920 21566 31096
rect 21790 30920 21824 31096
rect 22048 30920 22082 31096
rect 22306 30920 22340 31096
rect 22564 30920 22598 31096
rect 22822 30920 22856 31096
rect 23080 30920 23114 31096
rect 23338 30920 23372 31096
rect 20304 30827 20472 30861
rect 20562 30827 20730 30861
rect 20820 30827 20988 30861
rect 21078 30827 21246 30861
rect 21336 30827 21504 30861
rect 21594 30827 21762 30861
rect 21852 30827 22020 30861
rect 22110 30827 22278 30861
rect 22368 30827 22536 30861
rect 22626 30827 22794 30861
rect 22884 30827 23052 30861
rect 23142 30827 23310 30861
rect 20562 30719 20730 30753
rect 21336 30719 21504 30753
rect 21594 30719 21762 30753
rect 22368 30719 22536 30753
rect 22626 30719 22794 30753
rect 20242 30493 20276 30669
rect 20500 30493 20534 30669
rect 20758 30493 20792 30669
rect 21016 30493 21050 30669
rect 21274 30493 21308 30669
rect 21532 30493 21566 30669
rect 21790 30493 21824 30669
rect 22048 30493 22082 30669
rect 22306 30493 22340 30669
rect 22564 30493 22598 30669
rect 22822 30493 22856 30669
rect 23080 30493 23114 30669
rect 23338 30493 23372 30669
rect 20304 30409 20472 30443
rect 20820 30409 20988 30443
rect 21078 30409 21246 30443
rect 21852 30409 22020 30443
rect 22110 30409 22278 30443
rect 22884 30409 23052 30443
rect 23142 30409 23310 30443
rect 20304 30283 20472 30317
rect 20562 30283 20730 30317
rect 20820 30283 20988 30317
rect 21078 30283 21246 30317
rect 21336 30283 21504 30317
rect 21594 30283 21762 30317
rect 21852 30283 22020 30317
rect 22110 30283 22278 30317
rect 22368 30283 22536 30317
rect 22626 30283 22794 30317
rect 22884 30283 23052 30317
rect 23142 30283 23310 30317
rect 20242 30173 20276 30233
rect 20500 30173 20534 30233
rect 20758 30173 20792 30233
rect 21016 30173 21050 30233
rect 21274 30173 21308 30233
rect 21532 30173 21566 30233
rect 21790 30173 21824 30233
rect 22048 30173 22082 30233
rect 22306 30173 22340 30233
rect 22564 30173 22598 30233
rect 22822 30173 22856 30233
rect 23080 30173 23114 30233
rect 23338 30173 23372 30233
rect 19708 30096 20108 30106
rect 19708 30026 20076 30096
rect 20076 30026 20108 30096
rect 19708 30016 20108 30026
rect 20278 29996 23328 30046
rect 23678 31546 23718 31566
rect 23678 29656 23718 31546
rect 23678 29626 23718 29656
rect 18728 29586 18788 29626
rect 18788 29586 23648 29626
rect 23648 29586 23718 29626
rect 23948 31866 23988 31896
rect 23948 29316 23988 31866
rect 23948 29296 23988 29316
rect 18468 29256 18548 29296
rect 18548 29256 23918 29296
rect 23918 29256 23988 29296
rect 24388 31196 24508 31596
rect 24188 29616 24244 30056
rect 24244 29616 24278 30056
rect 24278 29616 24288 30056
rect 22288 29050 23408 29056
rect 12603 28963 12637 28997
rect 12695 28963 12729 28997
rect 12787 28963 12821 28997
rect 12879 28963 12913 28997
rect 12971 28963 13005 28997
rect 13063 28963 13097 28997
rect 13155 28963 13189 28997
rect 13247 28963 13281 28997
rect 13339 28963 13373 28997
rect 13431 28963 13465 28997
rect 13523 28963 13557 28997
rect 22288 29016 22340 29050
rect 22340 29016 23408 29050
rect 22288 28976 23408 29016
rect 22392 28798 22789 28904
rect 23591 28798 23988 28904
rect 24390 28800 24496 29197
rect 25625 31625 25659 31801
rect 25883 31625 25917 31801
rect 26141 31625 26175 31801
rect 25687 31541 25855 31575
rect 25945 31541 26113 31575
rect 26408 31636 26508 31816
rect 25687 30896 25855 30930
rect 25945 30896 26113 30930
rect 25625 30661 25659 30837
rect 25883 30661 25917 30837
rect 26141 30661 26175 30837
rect 26408 30656 26508 30836
rect 25625 30165 25659 30341
rect 25883 30165 25917 30341
rect 26141 30165 26175 30341
rect 25687 30081 25855 30115
rect 25945 30081 26113 30115
rect 26408 30176 26508 30356
rect 25335 29431 25369 29465
rect 25427 29431 25461 29465
rect 25519 29431 25553 29465
rect 25611 29431 25645 29465
rect 25703 29431 25737 29465
rect 25795 29431 25829 29465
rect 25887 29431 25921 29465
rect 25979 29431 26013 29465
rect 26071 29431 26105 29465
rect 26163 29431 26197 29465
rect 26255 29431 26289 29465
rect 25450 29153 25938 29160
rect 25450 29126 25458 29153
rect 25458 29126 25492 29153
rect 25492 29126 25542 29153
rect 25542 29126 25576 29153
rect 25576 29126 25626 29153
rect 25626 29126 25660 29153
rect 25660 29126 25710 29153
rect 25710 29126 25744 29153
rect 25744 29126 25794 29153
rect 25794 29126 25828 29153
rect 25828 29126 25878 29153
rect 25878 29126 25912 29153
rect 25912 29126 25938 29153
rect 26062 29060 26110 29224
rect 25335 28887 25369 28921
rect 25427 28887 25461 28921
rect 25519 28887 25553 28921
rect 25611 28887 25645 28921
rect 25703 28887 25737 28921
rect 25795 28887 25829 28921
rect 25887 28887 25921 28921
rect 25979 28887 26013 28921
rect 26071 28887 26105 28921
rect 26163 28887 26197 28921
rect 26255 28887 26289 28921
rect 13075 25728 13243 25762
rect 13333 25728 13501 25762
rect 13013 25493 13047 25669
rect 13271 25493 13305 25669
rect 13529 25493 13563 25669
rect 13796 25488 13896 25668
rect 5856 25268 5906 25308
rect 5906 25268 11306 25308
rect 11306 25268 11376 25308
rect 5856 25228 5896 25268
rect 5856 22698 5896 25228
rect 5856 22668 5896 22698
rect 6116 24938 6176 24978
rect 6176 24938 11026 24978
rect 11026 24938 11106 24978
rect 6116 24908 6156 24938
rect 6116 23038 6156 24908
rect 6116 22998 6156 23038
rect 7136 24568 7464 24608
rect 7464 24568 7706 24608
rect 7706 24568 10716 24608
rect 7630 24292 7664 24468
rect 7888 24292 7922 24468
rect 8146 24292 8180 24468
rect 8404 24292 8438 24468
rect 8662 24292 8696 24468
rect 8920 24292 8954 24468
rect 9178 24292 9212 24468
rect 9436 24292 9470 24468
rect 9694 24292 9728 24468
rect 9952 24292 9986 24468
rect 10210 24292 10244 24468
rect 10468 24292 10502 24468
rect 10726 24292 10760 24468
rect 7692 24199 7860 24233
rect 7950 24199 8118 24233
rect 8208 24199 8376 24233
rect 8466 24199 8634 24233
rect 8724 24199 8892 24233
rect 8982 24199 9150 24233
rect 9240 24199 9408 24233
rect 9498 24199 9666 24233
rect 9756 24199 9924 24233
rect 10014 24199 10182 24233
rect 10272 24199 10440 24233
rect 10530 24199 10698 24233
rect 7950 24091 8118 24125
rect 8724 24091 8892 24125
rect 8982 24091 9150 24125
rect 9756 24091 9924 24125
rect 10014 24091 10182 24125
rect 7630 23865 7664 24041
rect 7888 23865 7922 24041
rect 8146 23865 8180 24041
rect 8404 23865 8438 24041
rect 8662 23865 8696 24041
rect 8920 23865 8954 24041
rect 9178 23865 9212 24041
rect 9436 23865 9470 24041
rect 9694 23865 9728 24041
rect 9952 23865 9986 24041
rect 10210 23865 10244 24041
rect 10468 23865 10502 24041
rect 10726 23865 10760 24041
rect 7692 23781 7860 23815
rect 8208 23781 8376 23815
rect 8466 23781 8634 23815
rect 9240 23781 9408 23815
rect 9498 23781 9666 23815
rect 10272 23781 10440 23815
rect 10530 23781 10698 23815
rect 7692 23655 7860 23689
rect 7950 23655 8118 23689
rect 8208 23655 8376 23689
rect 8466 23655 8634 23689
rect 8724 23655 8892 23689
rect 8982 23655 9150 23689
rect 9240 23655 9408 23689
rect 9498 23655 9666 23689
rect 9756 23655 9924 23689
rect 10014 23655 10182 23689
rect 10272 23655 10440 23689
rect 10530 23655 10698 23689
rect 7630 23545 7664 23605
rect 7888 23545 7922 23605
rect 8146 23545 8180 23605
rect 8404 23545 8438 23605
rect 8662 23545 8696 23605
rect 8920 23545 8954 23605
rect 9178 23545 9212 23605
rect 9436 23545 9470 23605
rect 9694 23545 9728 23605
rect 9952 23545 9986 23605
rect 10210 23545 10244 23605
rect 10468 23545 10502 23605
rect 10726 23545 10760 23605
rect 7096 23468 7496 23478
rect 7096 23398 7464 23468
rect 7464 23398 7496 23468
rect 7096 23388 7496 23398
rect 7666 23368 10716 23418
rect 11066 24918 11106 24938
rect 11066 23028 11106 24918
rect 11066 22998 11106 23028
rect 6116 22958 6176 22998
rect 6176 22958 11036 22998
rect 11036 22958 11106 22998
rect 11336 25238 11376 25268
rect 11336 22688 11376 25238
rect 11336 22668 11376 22688
rect 5856 22628 5936 22668
rect 5936 22628 11306 22668
rect 11306 22628 11376 22668
rect 25783 25598 25951 25632
rect 26041 25598 26209 25632
rect 25721 25363 25755 25539
rect 25979 25363 26013 25539
rect 26237 25363 26271 25539
rect 11776 24568 11896 24968
rect 11576 22988 11632 23428
rect 11632 22988 11666 23428
rect 11666 22988 11676 23428
rect 9676 22422 10796 22428
rect 9676 22388 9728 22422
rect 9728 22388 10796 22422
rect 9676 22348 10796 22388
rect 9780 22170 10177 22276
rect 10979 22170 11376 22276
rect 11778 22172 11884 22569
rect 13013 24997 13047 25173
rect 13271 24997 13305 25173
rect 13529 24997 13563 25173
rect 13075 24913 13243 24947
rect 13333 24913 13501 24947
rect 26504 25358 26604 25538
rect 13796 25008 13896 25188
rect 13075 24268 13243 24302
rect 13333 24268 13501 24302
rect 13013 24033 13047 24209
rect 13271 24033 13305 24209
rect 13529 24033 13563 24209
rect 13796 24028 13896 24208
rect 13013 23537 13047 23713
rect 13271 23537 13305 23713
rect 13529 23537 13563 23713
rect 13075 23453 13243 23487
rect 13333 23453 13501 23487
rect 13796 23548 13896 23728
rect 12723 22803 12757 22837
rect 12815 22803 12849 22837
rect 12907 22803 12941 22837
rect 12999 22803 13033 22837
rect 13091 22803 13125 22837
rect 13183 22803 13217 22837
rect 13275 22803 13309 22837
rect 13367 22803 13401 22837
rect 13459 22803 13493 22837
rect 13551 22803 13585 22837
rect 13643 22803 13677 22837
rect 12838 22525 13326 22532
rect 12838 22498 12846 22525
rect 12846 22498 12880 22525
rect 12880 22498 12930 22525
rect 12930 22498 12964 22525
rect 12964 22498 13014 22525
rect 13014 22498 13048 22525
rect 13048 22498 13098 22525
rect 13098 22498 13132 22525
rect 13132 22498 13182 22525
rect 13182 22498 13216 22525
rect 13216 22498 13266 22525
rect 13266 22498 13300 22525
rect 13300 22498 13326 22525
rect 13450 22432 13498 22596
rect 18564 25138 18614 25178
rect 18614 25138 24014 25178
rect 24014 25138 24084 25178
rect 18564 25098 18604 25138
rect 18564 22568 18604 25098
rect 18564 22538 18604 22568
rect 18824 24808 18884 24848
rect 18884 24808 23734 24848
rect 23734 24808 23814 24848
rect 18824 24778 18864 24808
rect 18824 22908 18864 24778
rect 18824 22868 18864 22908
rect 19844 24438 20172 24478
rect 20172 24438 20414 24478
rect 20414 24438 23424 24478
rect 20338 24162 20372 24338
rect 20596 24162 20630 24338
rect 20854 24162 20888 24338
rect 21112 24162 21146 24338
rect 21370 24162 21404 24338
rect 21628 24162 21662 24338
rect 21886 24162 21920 24338
rect 22144 24162 22178 24338
rect 22402 24162 22436 24338
rect 22660 24162 22694 24338
rect 22918 24162 22952 24338
rect 23176 24162 23210 24338
rect 23434 24162 23468 24338
rect 20400 24069 20568 24103
rect 20658 24069 20826 24103
rect 20916 24069 21084 24103
rect 21174 24069 21342 24103
rect 21432 24069 21600 24103
rect 21690 24069 21858 24103
rect 21948 24069 22116 24103
rect 22206 24069 22374 24103
rect 22464 24069 22632 24103
rect 22722 24069 22890 24103
rect 22980 24069 23148 24103
rect 23238 24069 23406 24103
rect 20658 23961 20826 23995
rect 21432 23961 21600 23995
rect 21690 23961 21858 23995
rect 22464 23961 22632 23995
rect 22722 23961 22890 23995
rect 20338 23735 20372 23911
rect 20596 23735 20630 23911
rect 20854 23735 20888 23911
rect 21112 23735 21146 23911
rect 21370 23735 21404 23911
rect 21628 23735 21662 23911
rect 21886 23735 21920 23911
rect 22144 23735 22178 23911
rect 22402 23735 22436 23911
rect 22660 23735 22694 23911
rect 22918 23735 22952 23911
rect 23176 23735 23210 23911
rect 23434 23735 23468 23911
rect 20400 23651 20568 23685
rect 20916 23651 21084 23685
rect 21174 23651 21342 23685
rect 21948 23651 22116 23685
rect 22206 23651 22374 23685
rect 22980 23651 23148 23685
rect 23238 23651 23406 23685
rect 20400 23525 20568 23559
rect 20658 23525 20826 23559
rect 20916 23525 21084 23559
rect 21174 23525 21342 23559
rect 21432 23525 21600 23559
rect 21690 23525 21858 23559
rect 21948 23525 22116 23559
rect 22206 23525 22374 23559
rect 22464 23525 22632 23559
rect 22722 23525 22890 23559
rect 22980 23525 23148 23559
rect 23238 23525 23406 23559
rect 20338 23415 20372 23475
rect 20596 23415 20630 23475
rect 20854 23415 20888 23475
rect 21112 23415 21146 23475
rect 21370 23415 21404 23475
rect 21628 23415 21662 23475
rect 21886 23415 21920 23475
rect 22144 23415 22178 23475
rect 22402 23415 22436 23475
rect 22660 23415 22694 23475
rect 22918 23415 22952 23475
rect 23176 23415 23210 23475
rect 23434 23415 23468 23475
rect 19804 23338 20204 23348
rect 19804 23268 20172 23338
rect 20172 23268 20204 23338
rect 19804 23258 20204 23268
rect 20374 23238 23424 23288
rect 23774 24788 23814 24808
rect 23774 22898 23814 24788
rect 23774 22868 23814 22898
rect 18824 22828 18884 22868
rect 18884 22828 23744 22868
rect 23744 22828 23814 22868
rect 24044 25108 24084 25138
rect 24044 22558 24084 25108
rect 24044 22538 24084 22558
rect 18564 22498 18644 22538
rect 18644 22498 24014 22538
rect 24014 22498 24084 22538
rect 24484 24438 24604 24838
rect 24284 22858 24340 23298
rect 24340 22858 24374 23298
rect 24374 22858 24384 23298
rect 12723 22259 12757 22293
rect 12815 22259 12849 22293
rect 12907 22259 12941 22293
rect 12999 22259 13033 22293
rect 13091 22259 13125 22293
rect 13183 22259 13217 22293
rect 13275 22259 13309 22293
rect 13367 22259 13401 22293
rect 13459 22259 13493 22293
rect 13551 22259 13585 22293
rect 13643 22259 13677 22293
rect 22384 22292 23504 22298
rect 22384 22258 22436 22292
rect 22436 22258 23504 22292
rect 22384 22218 23504 22258
rect 22488 22040 22885 22146
rect 23687 22040 24084 22146
rect 24486 22042 24592 22439
rect 25721 24867 25755 25043
rect 25979 24867 26013 25043
rect 26237 24867 26271 25043
rect 25783 24783 25951 24817
rect 26041 24783 26209 24817
rect 26504 24878 26604 25058
rect 25783 24138 25951 24172
rect 26041 24138 26209 24172
rect 25721 23903 25755 24079
rect 25979 23903 26013 24079
rect 26237 23903 26271 24079
rect 26504 23898 26604 24078
rect 25721 23407 25755 23583
rect 25979 23407 26013 23583
rect 26237 23407 26271 23583
rect 25783 23323 25951 23357
rect 26041 23323 26209 23357
rect 26504 23418 26604 23598
rect 25431 22673 25465 22707
rect 25523 22673 25557 22707
rect 25615 22673 25649 22707
rect 25707 22673 25741 22707
rect 25799 22673 25833 22707
rect 25891 22673 25925 22707
rect 25983 22673 26017 22707
rect 26075 22673 26109 22707
rect 26167 22673 26201 22707
rect 26259 22673 26293 22707
rect 26351 22673 26385 22707
rect 25546 22395 26034 22402
rect 25546 22368 25554 22395
rect 25554 22368 25588 22395
rect 25588 22368 25638 22395
rect 25638 22368 25672 22395
rect 25672 22368 25722 22395
rect 25722 22368 25756 22395
rect 25756 22368 25806 22395
rect 25806 22368 25840 22395
rect 25840 22368 25890 22395
rect 25890 22368 25924 22395
rect 25924 22368 25974 22395
rect 25974 22368 26008 22395
rect 26008 22368 26034 22395
rect 26158 22302 26206 22466
rect 25431 22129 25465 22163
rect 25523 22129 25557 22163
rect 25615 22129 25649 22163
rect 25707 22129 25741 22163
rect 25799 22129 25833 22163
rect 25891 22129 25925 22163
rect 25983 22129 26017 22163
rect 26075 22129 26109 22163
rect 26167 22129 26201 22163
rect 26259 22129 26293 22163
rect 26351 22129 26385 22163
rect 12951 18682 13119 18716
rect 13209 18682 13377 18716
rect 12889 18447 12923 18623
rect 13147 18447 13181 18623
rect 13405 18447 13439 18623
rect 13672 18442 13772 18622
rect 5732 18222 5782 18262
rect 5782 18222 11182 18262
rect 11182 18222 11252 18262
rect 5732 18182 5772 18222
rect 5732 15652 5772 18182
rect 5732 15622 5772 15652
rect 5992 17892 6052 17932
rect 6052 17892 10902 17932
rect 10902 17892 10982 17932
rect 5992 17862 6032 17892
rect 5992 15992 6032 17862
rect 5992 15952 6032 15992
rect 7012 17522 7340 17562
rect 7340 17522 7582 17562
rect 7582 17522 10592 17562
rect 7506 17246 7540 17422
rect 7764 17246 7798 17422
rect 8022 17246 8056 17422
rect 8280 17246 8314 17422
rect 8538 17246 8572 17422
rect 8796 17246 8830 17422
rect 9054 17246 9088 17422
rect 9312 17246 9346 17422
rect 9570 17246 9604 17422
rect 9828 17246 9862 17422
rect 10086 17246 10120 17422
rect 10344 17246 10378 17422
rect 10602 17246 10636 17422
rect 7568 17153 7736 17187
rect 7826 17153 7994 17187
rect 8084 17153 8252 17187
rect 8342 17153 8510 17187
rect 8600 17153 8768 17187
rect 8858 17153 9026 17187
rect 9116 17153 9284 17187
rect 9374 17153 9542 17187
rect 9632 17153 9800 17187
rect 9890 17153 10058 17187
rect 10148 17153 10316 17187
rect 10406 17153 10574 17187
rect 7826 17045 7994 17079
rect 8600 17045 8768 17079
rect 8858 17045 9026 17079
rect 9632 17045 9800 17079
rect 9890 17045 10058 17079
rect 7506 16819 7540 16995
rect 7764 16819 7798 16995
rect 8022 16819 8056 16995
rect 8280 16819 8314 16995
rect 8538 16819 8572 16995
rect 8796 16819 8830 16995
rect 9054 16819 9088 16995
rect 9312 16819 9346 16995
rect 9570 16819 9604 16995
rect 9828 16819 9862 16995
rect 10086 16819 10120 16995
rect 10344 16819 10378 16995
rect 10602 16819 10636 16995
rect 7568 16735 7736 16769
rect 8084 16735 8252 16769
rect 8342 16735 8510 16769
rect 9116 16735 9284 16769
rect 9374 16735 9542 16769
rect 10148 16735 10316 16769
rect 10406 16735 10574 16769
rect 7568 16609 7736 16643
rect 7826 16609 7994 16643
rect 8084 16609 8252 16643
rect 8342 16609 8510 16643
rect 8600 16609 8768 16643
rect 8858 16609 9026 16643
rect 9116 16609 9284 16643
rect 9374 16609 9542 16643
rect 9632 16609 9800 16643
rect 9890 16609 10058 16643
rect 10148 16609 10316 16643
rect 10406 16609 10574 16643
rect 7506 16499 7540 16559
rect 7764 16499 7798 16559
rect 8022 16499 8056 16559
rect 8280 16499 8314 16559
rect 8538 16499 8572 16559
rect 8796 16499 8830 16559
rect 9054 16499 9088 16559
rect 9312 16499 9346 16559
rect 9570 16499 9604 16559
rect 9828 16499 9862 16559
rect 10086 16499 10120 16559
rect 10344 16499 10378 16559
rect 10602 16499 10636 16559
rect 6972 16422 7372 16432
rect 6972 16352 7340 16422
rect 7340 16352 7372 16422
rect 6972 16342 7372 16352
rect 7542 16322 10592 16372
rect 10942 17872 10982 17892
rect 10942 15982 10982 17872
rect 10942 15952 10982 15982
rect 5992 15912 6052 15952
rect 6052 15912 10912 15952
rect 10912 15912 10982 15952
rect 11212 18192 11252 18222
rect 11212 15642 11252 18192
rect 11212 15622 11252 15642
rect 5732 15582 5812 15622
rect 5812 15582 11182 15622
rect 11182 15582 11252 15622
rect 26133 18552 26301 18586
rect 26391 18552 26559 18586
rect 26071 18317 26105 18493
rect 26329 18317 26363 18493
rect 26587 18317 26621 18493
rect 11652 17522 11772 17922
rect 11452 15942 11508 16382
rect 11508 15942 11542 16382
rect 11542 15942 11552 16382
rect 9552 15376 10672 15382
rect 9552 15342 9604 15376
rect 9604 15342 10672 15376
rect 9552 15302 10672 15342
rect 9656 15124 10053 15230
rect 10855 15124 11252 15230
rect 11654 15126 11760 15523
rect 12889 17951 12923 18127
rect 13147 17951 13181 18127
rect 13405 17951 13439 18127
rect 12951 17867 13119 17901
rect 13209 17867 13377 17901
rect 26854 18312 26954 18492
rect 13672 17962 13772 18142
rect 12951 17222 13119 17256
rect 13209 17222 13377 17256
rect 12889 16987 12923 17163
rect 13147 16987 13181 17163
rect 13405 16987 13439 17163
rect 13672 16982 13772 17162
rect 12889 16491 12923 16667
rect 13147 16491 13181 16667
rect 13405 16491 13439 16667
rect 12951 16407 13119 16441
rect 13209 16407 13377 16441
rect 13672 16502 13772 16682
rect 12599 15757 12633 15791
rect 12691 15757 12725 15791
rect 12783 15757 12817 15791
rect 12875 15757 12909 15791
rect 12967 15757 13001 15791
rect 13059 15757 13093 15791
rect 13151 15757 13185 15791
rect 13243 15757 13277 15791
rect 13335 15757 13369 15791
rect 13427 15757 13461 15791
rect 13519 15757 13553 15791
rect 12714 15479 13202 15486
rect 12714 15452 12722 15479
rect 12722 15452 12756 15479
rect 12756 15452 12806 15479
rect 12806 15452 12840 15479
rect 12840 15452 12890 15479
rect 12890 15452 12924 15479
rect 12924 15452 12974 15479
rect 12974 15452 13008 15479
rect 13008 15452 13058 15479
rect 13058 15452 13092 15479
rect 13092 15452 13142 15479
rect 13142 15452 13176 15479
rect 13176 15452 13202 15479
rect 13326 15386 13374 15550
rect 18914 18092 18964 18132
rect 18964 18092 24364 18132
rect 24364 18092 24434 18132
rect 18914 18052 18954 18092
rect 18914 15522 18954 18052
rect 18914 15492 18954 15522
rect 19174 17762 19234 17802
rect 19234 17762 24084 17802
rect 24084 17762 24164 17802
rect 19174 17732 19214 17762
rect 19174 15862 19214 17732
rect 19174 15822 19214 15862
rect 20194 17392 20522 17432
rect 20522 17392 20764 17432
rect 20764 17392 23774 17432
rect 20688 17116 20722 17292
rect 20946 17116 20980 17292
rect 21204 17116 21238 17292
rect 21462 17116 21496 17292
rect 21720 17116 21754 17292
rect 21978 17116 22012 17292
rect 22236 17116 22270 17292
rect 22494 17116 22528 17292
rect 22752 17116 22786 17292
rect 23010 17116 23044 17292
rect 23268 17116 23302 17292
rect 23526 17116 23560 17292
rect 23784 17116 23818 17292
rect 20750 17023 20918 17057
rect 21008 17023 21176 17057
rect 21266 17023 21434 17057
rect 21524 17023 21692 17057
rect 21782 17023 21950 17057
rect 22040 17023 22208 17057
rect 22298 17023 22466 17057
rect 22556 17023 22724 17057
rect 22814 17023 22982 17057
rect 23072 17023 23240 17057
rect 23330 17023 23498 17057
rect 23588 17023 23756 17057
rect 21008 16915 21176 16949
rect 21782 16915 21950 16949
rect 22040 16915 22208 16949
rect 22814 16915 22982 16949
rect 23072 16915 23240 16949
rect 20688 16689 20722 16865
rect 20946 16689 20980 16865
rect 21204 16689 21238 16865
rect 21462 16689 21496 16865
rect 21720 16689 21754 16865
rect 21978 16689 22012 16865
rect 22236 16689 22270 16865
rect 22494 16689 22528 16865
rect 22752 16689 22786 16865
rect 23010 16689 23044 16865
rect 23268 16689 23302 16865
rect 23526 16689 23560 16865
rect 23784 16689 23818 16865
rect 20750 16605 20918 16639
rect 21266 16605 21434 16639
rect 21524 16605 21692 16639
rect 22298 16605 22466 16639
rect 22556 16605 22724 16639
rect 23330 16605 23498 16639
rect 23588 16605 23756 16639
rect 20750 16479 20918 16513
rect 21008 16479 21176 16513
rect 21266 16479 21434 16513
rect 21524 16479 21692 16513
rect 21782 16479 21950 16513
rect 22040 16479 22208 16513
rect 22298 16479 22466 16513
rect 22556 16479 22724 16513
rect 22814 16479 22982 16513
rect 23072 16479 23240 16513
rect 23330 16479 23498 16513
rect 23588 16479 23756 16513
rect 20688 16369 20722 16429
rect 20946 16369 20980 16429
rect 21204 16369 21238 16429
rect 21462 16369 21496 16429
rect 21720 16369 21754 16429
rect 21978 16369 22012 16429
rect 22236 16369 22270 16429
rect 22494 16369 22528 16429
rect 22752 16369 22786 16429
rect 23010 16369 23044 16429
rect 23268 16369 23302 16429
rect 23526 16369 23560 16429
rect 23784 16369 23818 16429
rect 20154 16292 20554 16302
rect 20154 16222 20522 16292
rect 20522 16222 20554 16292
rect 20154 16212 20554 16222
rect 20724 16192 23774 16242
rect 24124 17742 24164 17762
rect 24124 15852 24164 17742
rect 24124 15822 24164 15852
rect 19174 15782 19234 15822
rect 19234 15782 24094 15822
rect 24094 15782 24164 15822
rect 24394 18062 24434 18092
rect 24394 15512 24434 18062
rect 24394 15492 24434 15512
rect 18914 15452 18994 15492
rect 18994 15452 24364 15492
rect 24364 15452 24434 15492
rect 24834 17392 24954 17792
rect 24634 15812 24690 16252
rect 24690 15812 24724 16252
rect 24724 15812 24734 16252
rect 12599 15213 12633 15247
rect 12691 15213 12725 15247
rect 12783 15213 12817 15247
rect 12875 15213 12909 15247
rect 12967 15213 13001 15247
rect 13059 15213 13093 15247
rect 13151 15213 13185 15247
rect 13243 15213 13277 15247
rect 13335 15213 13369 15247
rect 13427 15213 13461 15247
rect 13519 15213 13553 15247
rect 22734 15246 23854 15252
rect 22734 15212 22786 15246
rect 22786 15212 23854 15246
rect 22734 15172 23854 15212
rect 22838 14994 23235 15100
rect 24037 14994 24434 15100
rect 24836 14996 24942 15393
rect 26071 17821 26105 17997
rect 26329 17821 26363 17997
rect 26587 17821 26621 17997
rect 26133 17737 26301 17771
rect 26391 17737 26559 17771
rect 26854 17832 26954 18012
rect 26133 17092 26301 17126
rect 26391 17092 26559 17126
rect 26071 16857 26105 17033
rect 26329 16857 26363 17033
rect 26587 16857 26621 17033
rect 26854 16852 26954 17032
rect 26071 16361 26105 16537
rect 26329 16361 26363 16537
rect 26587 16361 26621 16537
rect 26133 16277 26301 16311
rect 26391 16277 26559 16311
rect 26854 16372 26954 16552
rect 25781 15627 25815 15661
rect 25873 15627 25907 15661
rect 25965 15627 25999 15661
rect 26057 15627 26091 15661
rect 26149 15627 26183 15661
rect 26241 15627 26275 15661
rect 26333 15627 26367 15661
rect 26425 15627 26459 15661
rect 26517 15627 26551 15661
rect 26609 15627 26643 15661
rect 26701 15627 26735 15661
rect 25896 15349 26384 15356
rect 25896 15322 25904 15349
rect 25904 15322 25938 15349
rect 25938 15322 25988 15349
rect 25988 15322 26022 15349
rect 26022 15322 26072 15349
rect 26072 15322 26106 15349
rect 26106 15322 26156 15349
rect 26156 15322 26190 15349
rect 26190 15322 26240 15349
rect 26240 15322 26274 15349
rect 26274 15322 26324 15349
rect 26324 15322 26358 15349
rect 26358 15322 26384 15349
rect 26508 15256 26556 15420
rect 25781 15083 25815 15117
rect 25873 15083 25907 15117
rect 25965 15083 25999 15117
rect 26057 15083 26091 15117
rect 26149 15083 26183 15117
rect 26241 15083 26275 15117
rect 26333 15083 26367 15117
rect 26425 15083 26459 15117
rect 26517 15083 26551 15117
rect 26609 15083 26643 15117
rect 26701 15083 26735 15117
<< metal1 >>
rect 25704 38756 26164 38776
rect 12916 38638 13376 38658
rect 12916 38458 12936 38638
rect 13356 38458 13376 38638
rect 25704 38576 25724 38756
rect 26144 38576 26164 38756
rect 25704 38510 26164 38576
rect 25704 38476 25723 38510
rect 25891 38476 25981 38510
rect 26149 38476 26164 38510
rect 25711 38470 25903 38476
rect 25969 38470 26161 38476
rect 12916 38392 13376 38458
rect 26624 38436 27464 38476
rect 12916 38358 12935 38392
rect 13103 38358 13193 38392
rect 13361 38358 13376 38392
rect 25484 38417 25744 38436
rect 25484 38416 25661 38417
rect 25695 38416 25744 38417
rect 12923 38352 13115 38358
rect 13181 38352 13373 38358
rect 13836 38318 14676 38358
rect 12696 38299 12956 38318
rect 12696 38298 12873 38299
rect 12907 38298 12956 38299
rect 12696 38118 12716 38298
rect 12936 38118 12956 38298
rect 12696 38098 12956 38118
rect 13096 38299 13196 38318
rect 13096 38123 13131 38299
rect 13165 38123 13196 38299
rect 13096 38018 13196 38123
rect 13336 38299 13596 38318
rect 13336 38298 13389 38299
rect 13423 38298 13596 38299
rect 13336 38118 13356 38298
rect 13576 38118 13596 38298
rect 13336 38098 13596 38118
rect 13636 38298 14676 38318
rect 13636 38118 13656 38298
rect 13756 38118 14556 38298
rect 13636 38098 14556 38118
rect 13836 38078 14556 38098
rect 14636 38078 14676 38298
rect 25484 38236 25504 38416
rect 25724 38236 25744 38416
rect 25484 38216 25744 38236
rect 25884 38417 25984 38436
rect 25884 38241 25919 38417
rect 25953 38241 25984 38417
rect 25884 38136 25984 38241
rect 26124 38417 26384 38436
rect 26124 38416 26177 38417
rect 26211 38416 26384 38417
rect 26124 38236 26144 38416
rect 26364 38236 26384 38416
rect 26124 38216 26384 38236
rect 26424 38416 27464 38436
rect 26424 38236 26444 38416
rect 26544 38236 27344 38416
rect 26424 38216 27344 38236
rect 26624 38196 27344 38216
rect 27424 38196 27464 38416
rect 26624 38176 27464 38196
rect 13836 38058 14676 38078
rect 18404 38096 24104 38116
rect 18404 38056 20234 38096
rect 23444 38056 24104 38096
rect 5616 37978 11316 37998
rect 5616 37938 7446 37978
rect 10656 37938 11316 37978
rect 5616 35258 5716 37938
rect 5756 37818 7446 37898
rect 10656 37818 11196 37898
rect 5756 37798 11196 37818
rect 5756 35398 5816 37798
rect 5916 37608 11016 37698
rect 5916 35588 5976 37608
rect 6016 37498 10926 37568
rect 6016 35698 6116 37498
rect 6890 37258 10626 37278
rect 6890 37238 7446 37258
rect 6890 37198 6996 37238
rect 6890 37178 7446 37198
rect 10606 37178 10626 37258
rect 6890 37158 10626 37178
rect 7486 37110 7546 37158
rect 7484 37098 7546 37110
rect 7736 37108 7796 37118
rect 7484 36922 7490 37098
rect 7524 36922 7546 37098
rect 7484 36910 7546 36922
rect 7696 37098 7846 37108
rect 7696 36988 7748 37098
rect 7782 36988 7846 37098
rect 7696 36928 7706 36988
rect 7816 36928 7846 36988
rect 7696 36922 7748 36928
rect 7782 36922 7846 36928
rect 7696 36918 7846 36922
rect 7956 37098 8086 37158
rect 8258 37108 8304 37110
rect 7956 36922 8006 37098
rect 8040 36922 8086 37098
rect 7956 36918 8086 36922
rect 8216 37098 8346 37108
rect 8216 36988 8264 37098
rect 8298 36988 8346 37098
rect 8216 36928 8226 36988
rect 8336 36928 8346 36988
rect 8216 36922 8264 36928
rect 8298 36922 8346 36928
rect 8216 36918 8346 36922
rect 8476 37098 8606 37158
rect 8476 36922 8522 37098
rect 8556 36922 8606 37098
rect 8476 36918 8606 36922
rect 8726 37098 8856 37118
rect 8726 36988 8780 37098
rect 8814 36988 8856 37098
rect 7486 36869 7546 36910
rect 7736 36908 7846 36918
rect 8000 36910 8046 36918
rect 8258 36910 8304 36918
rect 8516 36910 8562 36918
rect 7796 36869 7846 36908
rect 8726 36878 8736 36988
rect 8846 36878 8856 36988
rect 8986 37098 9116 37158
rect 9290 37108 9336 37110
rect 8986 36922 9038 37098
rect 9072 36922 9116 37098
rect 8986 36918 9116 36922
rect 9246 37098 9376 37108
rect 9246 36998 9296 37098
rect 9330 36998 9376 37098
rect 9246 36928 9256 36998
rect 9366 36928 9376 36998
rect 9246 36922 9296 36928
rect 9330 36922 9376 36928
rect 9246 36918 9376 36922
rect 9506 37098 9636 37158
rect 9506 36922 9554 37098
rect 9588 36922 9636 37098
rect 9506 36918 9636 36922
rect 9766 37098 9896 37118
rect 9766 36998 9812 37098
rect 9846 36998 9896 37098
rect 9032 36910 9078 36918
rect 9290 36910 9336 36918
rect 9548 36910 9594 36918
rect 8726 36869 8856 36878
rect 9766 36878 9776 36998
rect 9886 36878 9896 36998
rect 10026 37098 10156 37158
rect 10586 37110 10626 37158
rect 10322 37108 10368 37110
rect 10026 36922 10070 37098
rect 10104 36922 10156 37098
rect 10026 36918 10156 36922
rect 10276 37098 10406 37108
rect 10276 36998 10328 37098
rect 10362 36998 10406 37098
rect 10276 36928 10286 36998
rect 10396 36928 10406 36998
rect 10276 36922 10328 36928
rect 10362 36922 10406 36928
rect 10276 36918 10406 36922
rect 10580 37098 10626 37110
rect 10580 36922 10586 37098
rect 10620 36922 10626 37098
rect 10064 36910 10110 36918
rect 10322 36910 10368 36918
rect 10580 36910 10626 36922
rect 10586 36878 10626 36910
rect 9766 36869 9896 36878
rect 7486 36868 7732 36869
rect 7486 36863 7736 36868
rect 7796 36863 7990 36869
rect 8056 36863 8248 36869
rect 8314 36863 8506 36869
rect 8572 36863 9022 36869
rect 9088 36863 9280 36869
rect 9346 36863 9538 36869
rect 9604 36863 10054 36869
rect 10120 36863 10312 36869
rect 10376 36863 10626 36878
rect 7486 36829 7552 36863
rect 7720 36829 7736 36863
rect 7794 36829 7810 36863
rect 7978 36829 8068 36863
rect 8236 36829 8326 36863
rect 8494 36829 8584 36863
rect 8752 36829 8842 36863
rect 9010 36829 9100 36863
rect 9268 36829 9358 36863
rect 9526 36829 9616 36863
rect 9784 36829 9874 36863
rect 10042 36829 10132 36863
rect 10300 36829 10316 36863
rect 10376 36829 10390 36863
rect 10558 36829 10626 36863
rect 7486 36828 7736 36829
rect 7796 36828 7990 36829
rect 7540 36823 7732 36828
rect 7798 36823 7990 36828
rect 8056 36823 8248 36829
rect 8314 36823 8506 36829
rect 8572 36823 8764 36829
rect 8830 36823 9022 36829
rect 9088 36823 9280 36829
rect 9346 36823 9538 36829
rect 9604 36823 9796 36829
rect 9862 36823 10054 36829
rect 10120 36823 10312 36829
rect 10376 36828 10626 36829
rect 10378 36823 10570 36828
rect 8076 36778 8186 36788
rect 7798 36755 7990 36761
rect 8076 36755 8086 36778
rect 7794 36721 7810 36755
rect 7978 36721 8086 36755
rect 7798 36715 7990 36721
rect 7486 36683 7536 36688
rect 7484 36671 7536 36683
rect 7742 36678 7788 36683
rect 7484 36495 7490 36671
rect 7524 36495 7536 36671
rect 7484 36483 7536 36495
rect 7696 36671 7826 36678
rect 7696 36668 7748 36671
rect 7782 36668 7826 36671
rect 7696 36608 7706 36668
rect 7816 36608 7826 36668
rect 7696 36495 7748 36608
rect 7782 36495 7826 36608
rect 8000 36671 8046 36683
rect 8000 36578 8006 36671
rect 7696 36488 7826 36495
rect 7956 36558 8006 36578
rect 8040 36578 8046 36671
rect 8076 36618 8086 36721
rect 8176 36755 8186 36778
rect 10146 36778 10246 36788
rect 8572 36755 8764 36761
rect 8830 36755 9022 36761
rect 9604 36755 9796 36761
rect 9862 36755 10054 36761
rect 8176 36721 8584 36755
rect 8752 36721 8842 36755
rect 9010 36721 9616 36755
rect 9784 36721 9874 36755
rect 10042 36721 10058 36755
rect 8176 36618 8186 36721
rect 8572 36715 8764 36721
rect 8830 36715 9022 36721
rect 9604 36715 9796 36721
rect 9862 36715 10054 36721
rect 8258 36678 8304 36683
rect 8516 36678 8562 36683
rect 8774 36678 8820 36683
rect 9032 36678 9078 36683
rect 9290 36678 9336 36683
rect 9548 36678 9594 36683
rect 9806 36678 9852 36683
rect 8076 36608 8186 36618
rect 8216 36671 8346 36678
rect 8216 36668 8264 36671
rect 8298 36668 8346 36671
rect 8216 36608 8226 36668
rect 8336 36608 8346 36668
rect 8040 36558 8086 36578
rect 7956 36498 7966 36558
rect 8076 36498 8086 36558
rect 7956 36495 8006 36498
rect 8040 36495 8086 36498
rect 7956 36488 8086 36495
rect 8216 36495 8264 36608
rect 8298 36495 8346 36608
rect 8216 36488 8346 36495
rect 8476 36671 8606 36678
rect 8476 36558 8522 36671
rect 8556 36558 8606 36671
rect 8476 36498 8486 36558
rect 8596 36498 8606 36558
rect 8476 36495 8522 36498
rect 8556 36495 8606 36498
rect 8476 36488 8606 36495
rect 8726 36671 8856 36678
rect 8726 36668 8780 36671
rect 8814 36668 8856 36671
rect 8726 36608 8736 36668
rect 8846 36608 8856 36668
rect 8726 36495 8780 36608
rect 8814 36495 8856 36608
rect 8726 36488 8856 36495
rect 8996 36671 9126 36678
rect 8996 36558 9038 36671
rect 9072 36558 9126 36671
rect 8996 36498 9006 36558
rect 9116 36498 9126 36558
rect 8996 36495 9038 36498
rect 9072 36495 9126 36498
rect 8996 36488 9126 36495
rect 9246 36671 9376 36678
rect 9246 36668 9296 36671
rect 9330 36668 9376 36671
rect 9246 36608 9256 36668
rect 9366 36608 9376 36668
rect 9246 36495 9296 36608
rect 9330 36495 9376 36608
rect 9246 36488 9376 36495
rect 9506 36671 9636 36678
rect 9506 36558 9554 36671
rect 9588 36558 9636 36671
rect 9506 36498 9516 36558
rect 9626 36498 9636 36558
rect 9506 36495 9554 36498
rect 9588 36495 9636 36498
rect 9506 36488 9636 36495
rect 9766 36671 9896 36678
rect 9766 36668 9812 36671
rect 9846 36668 9896 36671
rect 9766 36608 9776 36668
rect 9886 36608 9896 36668
rect 9766 36495 9812 36608
rect 9846 36495 9896 36608
rect 10064 36671 10110 36683
rect 10064 36568 10070 36671
rect 9766 36488 9896 36495
rect 10016 36558 10070 36568
rect 10104 36568 10110 36671
rect 10146 36628 10156 36778
rect 10236 36628 10246 36778
rect 10322 36678 10368 36683
rect 10146 36598 10246 36628
rect 10104 36558 10146 36568
rect 10016 36498 10026 36558
rect 10136 36498 10146 36558
rect 10016 36495 10070 36498
rect 10104 36495 10146 36498
rect 10016 36488 10146 36495
rect 7742 36483 7788 36488
rect 8000 36483 8046 36488
rect 8258 36483 8304 36488
rect 8516 36483 8562 36488
rect 8774 36483 8820 36488
rect 9032 36483 9078 36488
rect 9290 36483 9336 36488
rect 9548 36483 9594 36488
rect 9806 36483 9852 36488
rect 10064 36483 10110 36488
rect 7486 36478 7536 36483
rect 7486 36451 7556 36478
rect 10176 36451 10246 36598
rect 10276 36671 10406 36678
rect 10276 36668 10328 36671
rect 10362 36668 10406 36671
rect 10276 36608 10286 36668
rect 10396 36608 10406 36668
rect 10276 36495 10328 36608
rect 10362 36495 10406 36608
rect 10276 36488 10406 36495
rect 10576 36671 10626 36688
rect 10576 36495 10586 36671
rect 10620 36495 10626 36671
rect 10322 36483 10368 36488
rect 10576 36478 10626 36495
rect 10546 36451 10626 36478
rect 7486 36448 7732 36451
rect 7486 36445 7736 36448
rect 8056 36445 8248 36451
rect 8314 36445 8506 36451
rect 9088 36445 9280 36451
rect 9346 36445 9538 36451
rect 10120 36445 10312 36451
rect 10378 36448 10626 36451
rect 10366 36445 10626 36448
rect 7486 36411 7552 36445
rect 7720 36411 7736 36445
rect 8052 36411 8068 36445
rect 8236 36411 8326 36445
rect 8494 36411 9100 36445
rect 9268 36411 9358 36445
rect 9526 36411 10132 36445
rect 10300 36411 10316 36445
rect 10366 36411 10390 36445
rect 10558 36411 10626 36445
rect 7486 36348 7736 36411
rect 8056 36405 8248 36411
rect 8314 36405 8506 36411
rect 9088 36405 9280 36411
rect 9346 36405 9538 36411
rect 10120 36405 10312 36411
rect 7486 36319 8256 36348
rect 8936 36338 8946 36368
rect 7486 36285 7552 36319
rect 7720 36285 7810 36319
rect 7978 36285 8068 36319
rect 8236 36285 8256 36319
rect 7486 36268 8256 36285
rect 8306 36319 8946 36338
rect 9166 36338 9176 36368
rect 10366 36348 10626 36411
rect 9166 36319 9806 36338
rect 8306 36285 8326 36319
rect 8494 36285 8584 36319
rect 8752 36285 8842 36319
rect 9010 36285 9100 36308
rect 9268 36285 9358 36319
rect 9526 36285 9616 36319
rect 9784 36285 9806 36319
rect 8306 36278 9806 36285
rect 9856 36319 10626 36348
rect 9856 36285 9874 36319
rect 10042 36285 10132 36319
rect 10300 36285 10390 36319
rect 10558 36285 10626 36319
rect 8936 36268 9176 36278
rect 7486 36248 8276 36268
rect 7486 36247 8300 36248
rect 7484 36235 8304 36247
rect 7484 36175 7490 36235
rect 7524 36175 7748 36235
rect 7782 36175 8006 36235
rect 8040 36175 8264 36235
rect 8298 36175 8304 36235
rect 7484 36163 8304 36175
rect 8496 36173 8511 36248
rect 8566 36173 8586 36248
rect 8496 36163 8586 36173
rect 8726 36235 8866 36248
rect 8726 36175 8780 36235
rect 8814 36175 8866 36235
rect 6890 36128 7376 36138
rect 6890 36008 6946 36128
rect 7366 36008 7376 36128
rect 6890 35998 7376 36008
rect 7486 36078 8300 36163
rect 8726 36078 8866 36175
rect 9011 36235 9101 36268
rect 9856 36248 10626 36285
rect 9011 36175 9038 36235
rect 9072 36175 9101 36235
rect 9011 36158 9101 36175
rect 9246 36235 9386 36248
rect 9246 36175 9296 36235
rect 9330 36175 9386 36235
rect 9246 36078 9386 36175
rect 9531 36173 9541 36248
rect 9596 36173 9606 36248
rect 9531 36163 9606 36173
rect 9806 36235 10626 36248
rect 9806 36175 9812 36235
rect 9846 36175 10070 36235
rect 10104 36175 10328 36235
rect 10362 36175 10586 36235
rect 10620 36175 10626 36235
rect 9806 36078 10626 36175
rect 7486 36058 10626 36078
rect 7486 35988 7506 36058
rect 10606 35988 10626 36058
rect 7486 35968 10626 35988
rect 10816 35698 10926 37498
rect 6016 35678 10926 35698
rect 6016 35628 7446 35678
rect 10656 35628 10926 35678
rect 10966 35588 11016 37608
rect 5916 35518 7446 35588
rect 10656 35518 11016 35588
rect 5916 35498 11016 35518
rect 11116 35398 11196 37798
rect 5756 35298 11196 35398
rect 11236 35258 11316 37938
rect 12836 37938 13456 38018
rect 12836 37838 12936 37938
rect 13356 37838 13456 37938
rect 13836 37838 14676 37878
rect 12696 37818 12956 37838
rect 11576 37658 11836 37678
rect 11576 37178 11596 37658
rect 11816 37178 11836 37658
rect 12696 37638 12716 37818
rect 12936 37638 12956 37818
rect 13336 37818 13596 37838
rect 12696 37627 12873 37638
rect 12907 37627 12956 37638
rect 12696 37618 12956 37627
rect 13125 37803 13171 37815
rect 13125 37627 13131 37803
rect 13165 37627 13171 37803
rect 12867 37615 12913 37618
rect 13125 37615 13171 37627
rect 13336 37638 13356 37818
rect 13576 37638 13596 37818
rect 13336 37627 13389 37638
rect 13423 37627 13596 37638
rect 13336 37618 13596 37627
rect 13636 37818 14376 37838
rect 13636 37638 13656 37818
rect 13756 37638 14376 37818
rect 13636 37618 14376 37638
rect 14456 37618 14676 37838
rect 13383 37615 13429 37618
rect 12923 37578 13115 37583
rect 13181 37578 13373 37583
rect 13836 37578 14676 37618
rect 12916 37577 13376 37578
rect 12916 37543 12935 37577
rect 13103 37543 13193 37577
rect 13361 37543 13376 37577
rect 12916 37478 13376 37543
rect 12916 37298 12936 37478
rect 13356 37298 13376 37478
rect 12916 37278 13376 37298
rect 11576 37158 11836 37178
rect 12916 37178 13376 37198
rect 12916 36998 12936 37178
rect 13356 36998 13376 37178
rect 12916 36932 13376 36998
rect 12916 36898 12935 36932
rect 13103 36898 13193 36932
rect 13361 36898 13376 36932
rect 12923 36892 13115 36898
rect 13181 36892 13373 36898
rect 13836 36858 14676 36898
rect 12696 36839 12956 36858
rect 12696 36838 12873 36839
rect 12907 36838 12956 36839
rect 12696 36658 12716 36838
rect 12936 36658 12956 36838
rect 12696 36638 12956 36658
rect 13096 36839 13196 36858
rect 13096 36663 13131 36839
rect 13165 36663 13196 36839
rect 13096 36558 13196 36663
rect 13336 36839 13596 36858
rect 13336 36838 13389 36839
rect 13423 36838 13596 36839
rect 13336 36658 13356 36838
rect 13576 36658 13596 36838
rect 13336 36638 13596 36658
rect 13636 36838 14676 36858
rect 13636 36658 13656 36838
rect 13756 36658 14556 36838
rect 13636 36638 14556 36658
rect 13836 36618 14556 36638
rect 14636 36618 14676 36838
rect 13836 36598 14676 36618
rect 12836 36478 13456 36558
rect 12836 36378 12936 36478
rect 13356 36378 13456 36478
rect 13836 36378 14676 36418
rect 12696 36358 12956 36378
rect 12696 36178 12716 36358
rect 12936 36178 12956 36358
rect 13336 36358 13596 36378
rect 12696 36167 12873 36178
rect 12907 36167 12956 36178
rect 12696 36158 12956 36167
rect 13125 36343 13171 36355
rect 13125 36167 13131 36343
rect 13165 36167 13171 36343
rect 12867 36155 12913 36158
rect 13125 36155 13171 36167
rect 13336 36178 13356 36358
rect 13576 36178 13596 36358
rect 13336 36167 13389 36178
rect 13423 36167 13596 36178
rect 13336 36158 13596 36167
rect 13636 36358 14376 36378
rect 13636 36178 13656 36358
rect 13756 36178 14376 36358
rect 13636 36158 14376 36178
rect 14456 36158 14676 36378
rect 13383 36155 13429 36158
rect 12923 36118 13115 36123
rect 13181 36118 13373 36123
rect 13836 36118 14676 36158
rect 12916 36117 13376 36118
rect 12916 36083 12935 36117
rect 13103 36083 13193 36117
rect 13361 36083 13376 36117
rect 12916 36018 13376 36083
rect 12916 35838 12936 36018
rect 13356 35838 13376 36018
rect 12916 35818 13376 35838
rect 12554 35478 13566 35498
rect 12554 35418 12576 35478
rect 13536 35467 13566 35478
rect 13537 35433 13566 35467
rect 13536 35418 13566 35433
rect 12554 35402 13566 35418
rect 18404 35376 18504 38056
rect 18544 37936 20234 38016
rect 23444 37936 23984 38016
rect 18544 37916 23984 37936
rect 18544 35516 18604 37916
rect 18704 37726 23804 37816
rect 18704 35706 18764 37726
rect 18804 37616 23714 37686
rect 18804 35816 18904 37616
rect 19678 37376 23414 37396
rect 19678 37356 20234 37376
rect 19678 37316 19784 37356
rect 19678 37296 20234 37316
rect 23394 37296 23414 37376
rect 19678 37276 23414 37296
rect 20274 37228 20334 37276
rect 20272 37216 20334 37228
rect 20524 37226 20584 37236
rect 20272 37040 20278 37216
rect 20312 37040 20334 37216
rect 20272 37028 20334 37040
rect 20484 37216 20634 37226
rect 20484 37106 20536 37216
rect 20570 37106 20634 37216
rect 20484 37046 20494 37106
rect 20604 37046 20634 37106
rect 20484 37040 20536 37046
rect 20570 37040 20634 37046
rect 20484 37036 20634 37040
rect 20744 37216 20874 37276
rect 21046 37226 21092 37228
rect 20744 37040 20794 37216
rect 20828 37040 20874 37216
rect 20744 37036 20874 37040
rect 21004 37216 21134 37226
rect 21004 37106 21052 37216
rect 21086 37106 21134 37216
rect 21004 37046 21014 37106
rect 21124 37046 21134 37106
rect 21004 37040 21052 37046
rect 21086 37040 21134 37046
rect 21004 37036 21134 37040
rect 21264 37216 21394 37276
rect 21264 37040 21310 37216
rect 21344 37040 21394 37216
rect 21264 37036 21394 37040
rect 21514 37216 21644 37236
rect 21514 37106 21568 37216
rect 21602 37106 21644 37216
rect 20274 36987 20334 37028
rect 20524 37026 20634 37036
rect 20788 37028 20834 37036
rect 21046 37028 21092 37036
rect 21304 37028 21350 37036
rect 20584 36987 20634 37026
rect 21514 36996 21524 37106
rect 21634 36996 21644 37106
rect 21774 37216 21904 37276
rect 22078 37226 22124 37228
rect 21774 37040 21826 37216
rect 21860 37040 21904 37216
rect 21774 37036 21904 37040
rect 22034 37216 22164 37226
rect 22034 37116 22084 37216
rect 22118 37116 22164 37216
rect 22034 37046 22044 37116
rect 22154 37046 22164 37116
rect 22034 37040 22084 37046
rect 22118 37040 22164 37046
rect 22034 37036 22164 37040
rect 22294 37216 22424 37276
rect 22294 37040 22342 37216
rect 22376 37040 22424 37216
rect 22294 37036 22424 37040
rect 22554 37216 22684 37236
rect 22554 37116 22600 37216
rect 22634 37116 22684 37216
rect 21820 37028 21866 37036
rect 22078 37028 22124 37036
rect 22336 37028 22382 37036
rect 21514 36987 21644 36996
rect 22554 36996 22564 37116
rect 22674 36996 22684 37116
rect 22814 37216 22944 37276
rect 23374 37228 23414 37276
rect 23110 37226 23156 37228
rect 22814 37040 22858 37216
rect 22892 37040 22944 37216
rect 22814 37036 22944 37040
rect 23064 37216 23194 37226
rect 23064 37116 23116 37216
rect 23150 37116 23194 37216
rect 23064 37046 23074 37116
rect 23184 37046 23194 37116
rect 23064 37040 23116 37046
rect 23150 37040 23194 37046
rect 23064 37036 23194 37040
rect 23368 37216 23414 37228
rect 23368 37040 23374 37216
rect 23408 37040 23414 37216
rect 22852 37028 22898 37036
rect 23110 37028 23156 37036
rect 23368 37028 23414 37040
rect 23374 36996 23414 37028
rect 22554 36987 22684 36996
rect 20274 36986 20520 36987
rect 20274 36981 20524 36986
rect 20584 36981 20778 36987
rect 20844 36981 21036 36987
rect 21102 36981 21294 36987
rect 21360 36981 21810 36987
rect 21876 36981 22068 36987
rect 22134 36981 22326 36987
rect 22392 36981 22842 36987
rect 22908 36981 23100 36987
rect 23164 36981 23414 36996
rect 20274 36947 20340 36981
rect 20508 36947 20524 36981
rect 20582 36947 20598 36981
rect 20766 36947 20856 36981
rect 21024 36947 21114 36981
rect 21282 36947 21372 36981
rect 21540 36947 21630 36981
rect 21798 36947 21888 36981
rect 22056 36947 22146 36981
rect 22314 36947 22404 36981
rect 22572 36947 22662 36981
rect 22830 36947 22920 36981
rect 23088 36947 23104 36981
rect 23164 36947 23178 36981
rect 23346 36947 23414 36981
rect 20274 36946 20524 36947
rect 20584 36946 20778 36947
rect 20328 36941 20520 36946
rect 20586 36941 20778 36946
rect 20844 36941 21036 36947
rect 21102 36941 21294 36947
rect 21360 36941 21552 36947
rect 21618 36941 21810 36947
rect 21876 36941 22068 36947
rect 22134 36941 22326 36947
rect 22392 36941 22584 36947
rect 22650 36941 22842 36947
rect 22908 36941 23100 36947
rect 23164 36946 23414 36947
rect 23166 36941 23358 36946
rect 20864 36896 20974 36906
rect 20586 36873 20778 36879
rect 20864 36873 20874 36896
rect 20582 36839 20598 36873
rect 20766 36839 20874 36873
rect 20586 36833 20778 36839
rect 20274 36801 20324 36806
rect 20272 36789 20324 36801
rect 20530 36796 20576 36801
rect 20272 36613 20278 36789
rect 20312 36613 20324 36789
rect 20272 36601 20324 36613
rect 20484 36789 20614 36796
rect 20484 36786 20536 36789
rect 20570 36786 20614 36789
rect 20484 36726 20494 36786
rect 20604 36726 20614 36786
rect 20484 36613 20536 36726
rect 20570 36613 20614 36726
rect 20788 36789 20834 36801
rect 20788 36696 20794 36789
rect 20484 36606 20614 36613
rect 20744 36676 20794 36696
rect 20828 36696 20834 36789
rect 20864 36736 20874 36839
rect 20964 36873 20974 36896
rect 22934 36896 23034 36906
rect 21360 36873 21552 36879
rect 21618 36873 21810 36879
rect 22392 36873 22584 36879
rect 22650 36873 22842 36879
rect 20964 36839 21372 36873
rect 21540 36839 21630 36873
rect 21798 36839 22404 36873
rect 22572 36839 22662 36873
rect 22830 36839 22846 36873
rect 20964 36736 20974 36839
rect 21360 36833 21552 36839
rect 21618 36833 21810 36839
rect 22392 36833 22584 36839
rect 22650 36833 22842 36839
rect 21046 36796 21092 36801
rect 21304 36796 21350 36801
rect 21562 36796 21608 36801
rect 21820 36796 21866 36801
rect 22078 36796 22124 36801
rect 22336 36796 22382 36801
rect 22594 36796 22640 36801
rect 20864 36726 20974 36736
rect 21004 36789 21134 36796
rect 21004 36786 21052 36789
rect 21086 36786 21134 36789
rect 21004 36726 21014 36786
rect 21124 36726 21134 36786
rect 20828 36676 20874 36696
rect 20744 36616 20754 36676
rect 20864 36616 20874 36676
rect 20744 36613 20794 36616
rect 20828 36613 20874 36616
rect 20744 36606 20874 36613
rect 21004 36613 21052 36726
rect 21086 36613 21134 36726
rect 21004 36606 21134 36613
rect 21264 36789 21394 36796
rect 21264 36676 21310 36789
rect 21344 36676 21394 36789
rect 21264 36616 21274 36676
rect 21384 36616 21394 36676
rect 21264 36613 21310 36616
rect 21344 36613 21394 36616
rect 21264 36606 21394 36613
rect 21514 36789 21644 36796
rect 21514 36786 21568 36789
rect 21602 36786 21644 36789
rect 21514 36726 21524 36786
rect 21634 36726 21644 36786
rect 21514 36613 21568 36726
rect 21602 36613 21644 36726
rect 21514 36606 21644 36613
rect 21784 36789 21914 36796
rect 21784 36676 21826 36789
rect 21860 36676 21914 36789
rect 21784 36616 21794 36676
rect 21904 36616 21914 36676
rect 21784 36613 21826 36616
rect 21860 36613 21914 36616
rect 21784 36606 21914 36613
rect 22034 36789 22164 36796
rect 22034 36786 22084 36789
rect 22118 36786 22164 36789
rect 22034 36726 22044 36786
rect 22154 36726 22164 36786
rect 22034 36613 22084 36726
rect 22118 36613 22164 36726
rect 22034 36606 22164 36613
rect 22294 36789 22424 36796
rect 22294 36676 22342 36789
rect 22376 36676 22424 36789
rect 22294 36616 22304 36676
rect 22414 36616 22424 36676
rect 22294 36613 22342 36616
rect 22376 36613 22424 36616
rect 22294 36606 22424 36613
rect 22554 36789 22684 36796
rect 22554 36786 22600 36789
rect 22634 36786 22684 36789
rect 22554 36726 22564 36786
rect 22674 36726 22684 36786
rect 22554 36613 22600 36726
rect 22634 36613 22684 36726
rect 22852 36789 22898 36801
rect 22852 36686 22858 36789
rect 22554 36606 22684 36613
rect 22804 36676 22858 36686
rect 22892 36686 22898 36789
rect 22934 36746 22944 36896
rect 23024 36746 23034 36896
rect 23110 36796 23156 36801
rect 22934 36716 23034 36746
rect 22892 36676 22934 36686
rect 22804 36616 22814 36676
rect 22924 36616 22934 36676
rect 22804 36613 22858 36616
rect 22892 36613 22934 36616
rect 22804 36606 22934 36613
rect 20530 36601 20576 36606
rect 20788 36601 20834 36606
rect 21046 36601 21092 36606
rect 21304 36601 21350 36606
rect 21562 36601 21608 36606
rect 21820 36601 21866 36606
rect 22078 36601 22124 36606
rect 22336 36601 22382 36606
rect 22594 36601 22640 36606
rect 22852 36601 22898 36606
rect 20274 36596 20324 36601
rect 20274 36569 20344 36596
rect 22964 36569 23034 36716
rect 23064 36789 23194 36796
rect 23064 36786 23116 36789
rect 23150 36786 23194 36789
rect 23064 36726 23074 36786
rect 23184 36726 23194 36786
rect 23064 36613 23116 36726
rect 23150 36613 23194 36726
rect 23064 36606 23194 36613
rect 23364 36789 23414 36806
rect 23364 36613 23374 36789
rect 23408 36613 23414 36789
rect 23110 36601 23156 36606
rect 23364 36596 23414 36613
rect 23334 36569 23414 36596
rect 20274 36566 20520 36569
rect 20274 36563 20524 36566
rect 20844 36563 21036 36569
rect 21102 36563 21294 36569
rect 21876 36563 22068 36569
rect 22134 36563 22326 36569
rect 22908 36563 23100 36569
rect 23166 36566 23414 36569
rect 23154 36563 23414 36566
rect 20274 36529 20340 36563
rect 20508 36529 20524 36563
rect 20840 36529 20856 36563
rect 21024 36529 21114 36563
rect 21282 36529 21888 36563
rect 22056 36529 22146 36563
rect 22314 36529 22920 36563
rect 23088 36529 23104 36563
rect 23154 36529 23178 36563
rect 23346 36529 23414 36563
rect 20274 36466 20524 36529
rect 20844 36523 21036 36529
rect 21102 36523 21294 36529
rect 21876 36523 22068 36529
rect 22134 36523 22326 36529
rect 22908 36523 23100 36529
rect 20274 36437 21044 36466
rect 21724 36456 21734 36486
rect 20274 36403 20340 36437
rect 20508 36403 20598 36437
rect 20766 36403 20856 36437
rect 21024 36403 21044 36437
rect 20274 36386 21044 36403
rect 21094 36437 21734 36456
rect 21954 36456 21964 36486
rect 23154 36466 23414 36529
rect 21954 36437 22594 36456
rect 21094 36403 21114 36437
rect 21282 36403 21372 36437
rect 21540 36403 21630 36437
rect 21798 36403 21888 36426
rect 22056 36403 22146 36437
rect 22314 36403 22404 36437
rect 22572 36403 22594 36437
rect 21094 36396 22594 36403
rect 22644 36437 23414 36466
rect 22644 36403 22662 36437
rect 22830 36403 22920 36437
rect 23088 36403 23178 36437
rect 23346 36403 23414 36437
rect 21724 36386 21964 36396
rect 20274 36366 21064 36386
rect 20274 36365 21088 36366
rect 20272 36353 21092 36365
rect 20272 36293 20278 36353
rect 20312 36293 20536 36353
rect 20570 36293 20794 36353
rect 20828 36293 21052 36353
rect 21086 36293 21092 36353
rect 20272 36281 21092 36293
rect 21284 36291 21299 36366
rect 21354 36291 21374 36366
rect 21284 36281 21374 36291
rect 21514 36353 21654 36366
rect 21514 36293 21568 36353
rect 21602 36293 21654 36353
rect 19678 36246 20164 36256
rect 19678 36126 19734 36246
rect 20154 36126 20164 36246
rect 19678 36116 20164 36126
rect 20274 36196 21088 36281
rect 21514 36196 21654 36293
rect 21799 36353 21889 36386
rect 22644 36366 23414 36403
rect 21799 36293 21826 36353
rect 21860 36293 21889 36353
rect 21799 36276 21889 36293
rect 22034 36353 22174 36366
rect 22034 36293 22084 36353
rect 22118 36293 22174 36353
rect 22034 36196 22174 36293
rect 22319 36291 22329 36366
rect 22384 36291 22394 36366
rect 22319 36281 22394 36291
rect 22594 36353 23414 36366
rect 22594 36293 22600 36353
rect 22634 36293 22858 36353
rect 22892 36293 23116 36353
rect 23150 36293 23374 36353
rect 23408 36293 23414 36353
rect 22594 36196 23414 36293
rect 20274 36176 23414 36196
rect 20274 36106 20294 36176
rect 23394 36106 23414 36176
rect 20274 36086 23414 36106
rect 23604 35816 23714 37616
rect 18804 35796 23714 35816
rect 18804 35746 20234 35796
rect 23444 35746 23714 35796
rect 23754 35706 23804 37726
rect 18704 35636 20234 35706
rect 23444 35636 23804 35706
rect 18704 35616 23804 35636
rect 23904 35516 23984 37916
rect 18544 35416 23984 35516
rect 24024 35376 24104 38056
rect 25624 38056 26244 38136
rect 25624 37956 25724 38056
rect 26144 37956 26244 38056
rect 26624 37956 27464 37996
rect 25484 37936 25744 37956
rect 24364 37776 24624 37796
rect 24364 37296 24384 37776
rect 24604 37296 24624 37776
rect 25484 37756 25504 37936
rect 25724 37756 25744 37936
rect 26124 37936 26384 37956
rect 25484 37745 25661 37756
rect 25695 37745 25744 37756
rect 25484 37736 25744 37745
rect 25913 37921 25959 37933
rect 25913 37745 25919 37921
rect 25953 37745 25959 37921
rect 25655 37733 25701 37736
rect 25913 37733 25959 37745
rect 26124 37756 26144 37936
rect 26364 37756 26384 37936
rect 26124 37745 26177 37756
rect 26211 37745 26384 37756
rect 26124 37736 26384 37745
rect 26424 37936 27164 37956
rect 26424 37756 26444 37936
rect 26544 37756 27164 37936
rect 26424 37736 27164 37756
rect 27244 37736 27464 37956
rect 26171 37733 26217 37736
rect 25711 37696 25903 37701
rect 25969 37696 26161 37701
rect 26624 37696 27464 37736
rect 25704 37695 26164 37696
rect 25704 37661 25723 37695
rect 25891 37661 25981 37695
rect 26149 37661 26164 37695
rect 25704 37596 26164 37661
rect 25704 37416 25724 37596
rect 26144 37416 26164 37596
rect 25704 37396 26164 37416
rect 24364 37276 24624 37296
rect 25704 37296 26164 37316
rect 25704 37116 25724 37296
rect 26144 37116 26164 37296
rect 25704 37050 26164 37116
rect 25704 37016 25723 37050
rect 25891 37016 25981 37050
rect 26149 37016 26164 37050
rect 25711 37010 25903 37016
rect 25969 37010 26161 37016
rect 26624 36976 27464 37016
rect 25484 36957 25744 36976
rect 25484 36956 25661 36957
rect 25695 36956 25744 36957
rect 25484 36776 25504 36956
rect 25724 36776 25744 36956
rect 25484 36756 25744 36776
rect 25884 36957 25984 36976
rect 25884 36781 25919 36957
rect 25953 36781 25984 36957
rect 25884 36676 25984 36781
rect 26124 36957 26384 36976
rect 26124 36956 26177 36957
rect 26211 36956 26384 36957
rect 26124 36776 26144 36956
rect 26364 36776 26384 36956
rect 26124 36756 26384 36776
rect 26424 36956 27464 36976
rect 26424 36776 26444 36956
rect 26544 36776 27344 36956
rect 26424 36756 27344 36776
rect 26624 36736 27344 36756
rect 27424 36736 27464 36956
rect 26624 36716 27464 36736
rect 25624 36596 26244 36676
rect 25624 36496 25724 36596
rect 26144 36496 26244 36596
rect 26624 36496 27464 36536
rect 25484 36476 25744 36496
rect 25484 36296 25504 36476
rect 25724 36296 25744 36476
rect 26124 36476 26384 36496
rect 25484 36285 25661 36296
rect 25695 36285 25744 36296
rect 25484 36276 25744 36285
rect 25913 36461 25959 36473
rect 25913 36285 25919 36461
rect 25953 36285 25959 36461
rect 25655 36273 25701 36276
rect 25913 36273 25959 36285
rect 26124 36296 26144 36476
rect 26364 36296 26384 36476
rect 26124 36285 26177 36296
rect 26211 36285 26384 36296
rect 26124 36276 26384 36285
rect 26424 36476 27164 36496
rect 26424 36296 26444 36476
rect 26544 36296 27164 36476
rect 26424 36276 27164 36296
rect 27244 36276 27464 36496
rect 26171 36273 26217 36276
rect 25711 36236 25903 36241
rect 25969 36236 26161 36241
rect 26624 36236 27464 36276
rect 25704 36235 26164 36236
rect 25704 36201 25723 36235
rect 25891 36201 25981 36235
rect 26149 36201 26164 36235
rect 24204 36176 24344 36196
rect 24204 35736 24224 36176
rect 24324 35736 24344 36176
rect 25704 36136 26164 36201
rect 25704 35956 25724 36136
rect 26144 35956 26164 36136
rect 25704 35936 26164 35956
rect 24204 35716 24344 35736
rect 25342 35596 26354 35616
rect 25342 35536 25364 35596
rect 26324 35585 26354 35596
rect 26325 35551 26354 35585
rect 26324 35536 26354 35551
rect 25342 35520 26354 35536
rect 18404 35316 24104 35376
rect 24984 35356 25984 35376
rect 24384 35317 24584 35336
rect 24384 35316 24426 35317
rect 24532 35316 24584 35317
rect 5616 35198 11316 35258
rect 12196 35238 13196 35258
rect 12196 35058 12216 35238
rect 12396 35162 13196 35238
rect 12396 35128 12698 35162
rect 13186 35128 13196 35162
rect 12396 35058 13196 35128
rect 12196 35038 13196 35058
rect 13296 35238 13696 35258
rect 13296 35226 13496 35238
rect 13296 35062 13310 35226
rect 13358 35062 13496 35226
rect 13296 35058 13496 35062
rect 13676 35058 13696 35238
rect 22304 35194 23464 35196
rect 13296 35038 13696 35058
rect 22300 35176 23464 35194
rect 22300 35096 22324 35176
rect 23444 35096 23464 35176
rect 22300 35076 23464 35096
rect 22300 35024 22888 35076
rect 24384 35056 24404 35316
rect 12554 34938 13566 34954
rect 12554 34878 12576 34938
rect 13556 34878 13566 34938
rect 22300 34918 22428 35024
rect 22825 34918 22888 35024
rect 22300 34882 22888 34918
rect 23604 35036 24404 35056
rect 12554 34858 13566 34878
rect 23604 34856 23624 35036
rect 24564 34856 24584 35316
rect 24984 35176 25004 35356
rect 25184 35280 25984 35356
rect 25184 35246 25486 35280
rect 25974 35246 25984 35280
rect 25184 35176 25984 35246
rect 24984 35156 25984 35176
rect 26084 35356 26484 35376
rect 26084 35344 26284 35356
rect 26084 35180 26098 35344
rect 26146 35180 26284 35344
rect 26084 35176 26284 35180
rect 26464 35176 26484 35356
rect 26084 35156 26484 35176
rect 25342 35056 26354 35072
rect 25342 34996 25364 35056
rect 26344 34996 26354 35056
rect 25342 34976 26354 34996
rect 23604 34836 24584 34856
rect 12936 32712 13396 32732
rect 12936 32532 12956 32712
rect 13376 32532 13396 32712
rect 12936 32466 13396 32532
rect 12936 32432 12955 32466
rect 13123 32432 13213 32466
rect 13381 32432 13396 32466
rect 25668 32636 26128 32656
rect 25668 32456 25688 32636
rect 26108 32456 26128 32636
rect 12943 32426 13135 32432
rect 13201 32426 13393 32432
rect 13856 32392 14696 32432
rect 12716 32373 12976 32392
rect 12716 32372 12893 32373
rect 12927 32372 12976 32373
rect 12716 32192 12736 32372
rect 12956 32192 12976 32372
rect 12716 32172 12976 32192
rect 13116 32373 13216 32392
rect 13116 32197 13151 32373
rect 13185 32197 13216 32373
rect 13116 32092 13216 32197
rect 13356 32373 13616 32392
rect 13356 32372 13409 32373
rect 13443 32372 13616 32373
rect 13356 32192 13376 32372
rect 13596 32192 13616 32372
rect 13356 32172 13616 32192
rect 13656 32372 14696 32392
rect 13656 32192 13676 32372
rect 13776 32192 14576 32372
rect 13656 32172 14576 32192
rect 13856 32152 14576 32172
rect 14656 32152 14696 32372
rect 25668 32390 26128 32456
rect 25668 32356 25687 32390
rect 25855 32356 25945 32390
rect 26113 32356 26128 32390
rect 25675 32350 25867 32356
rect 25933 32350 26125 32356
rect 26588 32316 27428 32356
rect 13856 32132 14696 32152
rect 25448 32297 25708 32316
rect 25448 32296 25625 32297
rect 25659 32296 25708 32297
rect 25448 32116 25468 32296
rect 25688 32116 25708 32296
rect 25448 32096 25708 32116
rect 25848 32297 25948 32316
rect 25848 32121 25883 32297
rect 25917 32121 25948 32297
rect 5636 32052 11336 32072
rect 5636 32012 7466 32052
rect 10676 32012 11336 32052
rect 5636 29332 5736 32012
rect 5776 31892 7466 31972
rect 10676 31892 11216 31972
rect 5776 31872 11216 31892
rect 5776 29472 5836 31872
rect 5936 31682 11036 31772
rect 5936 29662 5996 31682
rect 6036 31572 10946 31642
rect 6036 29772 6136 31572
rect 6910 31332 10646 31352
rect 6910 31312 7466 31332
rect 6910 31272 7016 31312
rect 6910 31252 7466 31272
rect 10626 31252 10646 31332
rect 6910 31232 10646 31252
rect 7506 31184 7566 31232
rect 7504 31172 7566 31184
rect 7756 31182 7816 31192
rect 7504 30996 7510 31172
rect 7544 30996 7566 31172
rect 7504 30984 7566 30996
rect 7716 31172 7866 31182
rect 7716 31062 7768 31172
rect 7802 31062 7866 31172
rect 7716 31002 7726 31062
rect 7836 31002 7866 31062
rect 7716 30996 7768 31002
rect 7802 30996 7866 31002
rect 7716 30992 7866 30996
rect 7976 31172 8106 31232
rect 8278 31182 8324 31184
rect 7976 30996 8026 31172
rect 8060 30996 8106 31172
rect 7976 30992 8106 30996
rect 8236 31172 8366 31182
rect 8236 31062 8284 31172
rect 8318 31062 8366 31172
rect 8236 31002 8246 31062
rect 8356 31002 8366 31062
rect 8236 30996 8284 31002
rect 8318 30996 8366 31002
rect 8236 30992 8366 30996
rect 8496 31172 8626 31232
rect 8496 30996 8542 31172
rect 8576 30996 8626 31172
rect 8496 30992 8626 30996
rect 8746 31172 8876 31192
rect 8746 31062 8800 31172
rect 8834 31062 8876 31172
rect 7506 30943 7566 30984
rect 7756 30982 7866 30992
rect 8020 30984 8066 30992
rect 8278 30984 8324 30992
rect 8536 30984 8582 30992
rect 7816 30943 7866 30982
rect 8746 30952 8756 31062
rect 8866 30952 8876 31062
rect 9006 31172 9136 31232
rect 9310 31182 9356 31184
rect 9006 30996 9058 31172
rect 9092 30996 9136 31172
rect 9006 30992 9136 30996
rect 9266 31172 9396 31182
rect 9266 31072 9316 31172
rect 9350 31072 9396 31172
rect 9266 31002 9276 31072
rect 9386 31002 9396 31072
rect 9266 30996 9316 31002
rect 9350 30996 9396 31002
rect 9266 30992 9396 30996
rect 9526 31172 9656 31232
rect 9526 30996 9574 31172
rect 9608 30996 9656 31172
rect 9526 30992 9656 30996
rect 9786 31172 9916 31192
rect 9786 31072 9832 31172
rect 9866 31072 9916 31172
rect 9052 30984 9098 30992
rect 9310 30984 9356 30992
rect 9568 30984 9614 30992
rect 8746 30943 8876 30952
rect 9786 30952 9796 31072
rect 9906 30952 9916 31072
rect 10046 31172 10176 31232
rect 10606 31184 10646 31232
rect 10342 31182 10388 31184
rect 10046 30996 10090 31172
rect 10124 30996 10176 31172
rect 10046 30992 10176 30996
rect 10296 31172 10426 31182
rect 10296 31072 10348 31172
rect 10382 31072 10426 31172
rect 10296 31002 10306 31072
rect 10416 31002 10426 31072
rect 10296 30996 10348 31002
rect 10382 30996 10426 31002
rect 10296 30992 10426 30996
rect 10600 31172 10646 31184
rect 10600 30996 10606 31172
rect 10640 30996 10646 31172
rect 10084 30984 10130 30992
rect 10342 30984 10388 30992
rect 10600 30984 10646 30996
rect 10606 30952 10646 30984
rect 9786 30943 9916 30952
rect 7506 30942 7752 30943
rect 7506 30937 7756 30942
rect 7816 30937 8010 30943
rect 8076 30937 8268 30943
rect 8334 30937 8526 30943
rect 8592 30937 9042 30943
rect 9108 30937 9300 30943
rect 9366 30937 9558 30943
rect 9624 30937 10074 30943
rect 10140 30937 10332 30943
rect 10396 30937 10646 30952
rect 7506 30903 7572 30937
rect 7740 30903 7756 30937
rect 7814 30903 7830 30937
rect 7998 30903 8088 30937
rect 8256 30903 8346 30937
rect 8514 30903 8604 30937
rect 8772 30903 8862 30937
rect 9030 30903 9120 30937
rect 9288 30903 9378 30937
rect 9546 30903 9636 30937
rect 9804 30903 9894 30937
rect 10062 30903 10152 30937
rect 10320 30903 10336 30937
rect 10396 30903 10410 30937
rect 10578 30903 10646 30937
rect 7506 30902 7756 30903
rect 7816 30902 8010 30903
rect 7560 30897 7752 30902
rect 7818 30897 8010 30902
rect 8076 30897 8268 30903
rect 8334 30897 8526 30903
rect 8592 30897 8784 30903
rect 8850 30897 9042 30903
rect 9108 30897 9300 30903
rect 9366 30897 9558 30903
rect 9624 30897 9816 30903
rect 9882 30897 10074 30903
rect 10140 30897 10332 30903
rect 10396 30902 10646 30903
rect 10398 30897 10590 30902
rect 8096 30852 8206 30862
rect 7818 30829 8010 30835
rect 8096 30829 8106 30852
rect 7814 30795 7830 30829
rect 7998 30795 8106 30829
rect 7818 30789 8010 30795
rect 7506 30757 7556 30762
rect 7504 30745 7556 30757
rect 7762 30752 7808 30757
rect 7504 30569 7510 30745
rect 7544 30569 7556 30745
rect 7504 30557 7556 30569
rect 7716 30745 7846 30752
rect 7716 30742 7768 30745
rect 7802 30742 7846 30745
rect 7716 30682 7726 30742
rect 7836 30682 7846 30742
rect 7716 30569 7768 30682
rect 7802 30569 7846 30682
rect 8020 30745 8066 30757
rect 8020 30652 8026 30745
rect 7716 30562 7846 30569
rect 7976 30632 8026 30652
rect 8060 30652 8066 30745
rect 8096 30692 8106 30795
rect 8196 30829 8206 30852
rect 10166 30852 10266 30862
rect 8592 30829 8784 30835
rect 8850 30829 9042 30835
rect 9624 30829 9816 30835
rect 9882 30829 10074 30835
rect 8196 30795 8604 30829
rect 8772 30795 8862 30829
rect 9030 30795 9636 30829
rect 9804 30795 9894 30829
rect 10062 30795 10078 30829
rect 8196 30692 8206 30795
rect 8592 30789 8784 30795
rect 8850 30789 9042 30795
rect 9624 30789 9816 30795
rect 9882 30789 10074 30795
rect 8278 30752 8324 30757
rect 8536 30752 8582 30757
rect 8794 30752 8840 30757
rect 9052 30752 9098 30757
rect 9310 30752 9356 30757
rect 9568 30752 9614 30757
rect 9826 30752 9872 30757
rect 8096 30682 8206 30692
rect 8236 30745 8366 30752
rect 8236 30742 8284 30745
rect 8318 30742 8366 30745
rect 8236 30682 8246 30742
rect 8356 30682 8366 30742
rect 8060 30632 8106 30652
rect 7976 30572 7986 30632
rect 8096 30572 8106 30632
rect 7976 30569 8026 30572
rect 8060 30569 8106 30572
rect 7976 30562 8106 30569
rect 8236 30569 8284 30682
rect 8318 30569 8366 30682
rect 8236 30562 8366 30569
rect 8496 30745 8626 30752
rect 8496 30632 8542 30745
rect 8576 30632 8626 30745
rect 8496 30572 8506 30632
rect 8616 30572 8626 30632
rect 8496 30569 8542 30572
rect 8576 30569 8626 30572
rect 8496 30562 8626 30569
rect 8746 30745 8876 30752
rect 8746 30742 8800 30745
rect 8834 30742 8876 30745
rect 8746 30682 8756 30742
rect 8866 30682 8876 30742
rect 8746 30569 8800 30682
rect 8834 30569 8876 30682
rect 8746 30562 8876 30569
rect 9016 30745 9146 30752
rect 9016 30632 9058 30745
rect 9092 30632 9146 30745
rect 9016 30572 9026 30632
rect 9136 30572 9146 30632
rect 9016 30569 9058 30572
rect 9092 30569 9146 30572
rect 9016 30562 9146 30569
rect 9266 30745 9396 30752
rect 9266 30742 9316 30745
rect 9350 30742 9396 30745
rect 9266 30682 9276 30742
rect 9386 30682 9396 30742
rect 9266 30569 9316 30682
rect 9350 30569 9396 30682
rect 9266 30562 9396 30569
rect 9526 30745 9656 30752
rect 9526 30632 9574 30745
rect 9608 30632 9656 30745
rect 9526 30572 9536 30632
rect 9646 30572 9656 30632
rect 9526 30569 9574 30572
rect 9608 30569 9656 30572
rect 9526 30562 9656 30569
rect 9786 30745 9916 30752
rect 9786 30742 9832 30745
rect 9866 30742 9916 30745
rect 9786 30682 9796 30742
rect 9906 30682 9916 30742
rect 9786 30569 9832 30682
rect 9866 30569 9916 30682
rect 10084 30745 10130 30757
rect 10084 30642 10090 30745
rect 9786 30562 9916 30569
rect 10036 30632 10090 30642
rect 10124 30642 10130 30745
rect 10166 30702 10176 30852
rect 10256 30702 10266 30852
rect 10342 30752 10388 30757
rect 10166 30672 10266 30702
rect 10124 30632 10166 30642
rect 10036 30572 10046 30632
rect 10156 30572 10166 30632
rect 10036 30569 10090 30572
rect 10124 30569 10166 30572
rect 10036 30562 10166 30569
rect 7762 30557 7808 30562
rect 8020 30557 8066 30562
rect 8278 30557 8324 30562
rect 8536 30557 8582 30562
rect 8794 30557 8840 30562
rect 9052 30557 9098 30562
rect 9310 30557 9356 30562
rect 9568 30557 9614 30562
rect 9826 30557 9872 30562
rect 10084 30557 10130 30562
rect 7506 30552 7556 30557
rect 7506 30525 7576 30552
rect 10196 30525 10266 30672
rect 10296 30745 10426 30752
rect 10296 30742 10348 30745
rect 10382 30742 10426 30745
rect 10296 30682 10306 30742
rect 10416 30682 10426 30742
rect 10296 30569 10348 30682
rect 10382 30569 10426 30682
rect 10296 30562 10426 30569
rect 10596 30745 10646 30762
rect 10596 30569 10606 30745
rect 10640 30569 10646 30745
rect 10342 30557 10388 30562
rect 10596 30552 10646 30569
rect 10566 30525 10646 30552
rect 7506 30522 7752 30525
rect 7506 30519 7756 30522
rect 8076 30519 8268 30525
rect 8334 30519 8526 30525
rect 9108 30519 9300 30525
rect 9366 30519 9558 30525
rect 10140 30519 10332 30525
rect 10398 30522 10646 30525
rect 10386 30519 10646 30522
rect 7506 30485 7572 30519
rect 7740 30485 7756 30519
rect 8072 30485 8088 30519
rect 8256 30485 8346 30519
rect 8514 30485 9120 30519
rect 9288 30485 9378 30519
rect 9546 30485 10152 30519
rect 10320 30485 10336 30519
rect 10386 30485 10410 30519
rect 10578 30485 10646 30519
rect 7506 30422 7756 30485
rect 8076 30479 8268 30485
rect 8334 30479 8526 30485
rect 9108 30479 9300 30485
rect 9366 30479 9558 30485
rect 10140 30479 10332 30485
rect 7506 30393 8276 30422
rect 8956 30412 8966 30442
rect 7506 30359 7572 30393
rect 7740 30359 7830 30393
rect 7998 30359 8088 30393
rect 8256 30359 8276 30393
rect 7506 30342 8276 30359
rect 8326 30393 8966 30412
rect 9186 30412 9196 30442
rect 10386 30422 10646 30485
rect 9186 30393 9826 30412
rect 8326 30359 8346 30393
rect 8514 30359 8604 30393
rect 8772 30359 8862 30393
rect 9030 30359 9120 30382
rect 9288 30359 9378 30393
rect 9546 30359 9636 30393
rect 9804 30359 9826 30393
rect 8326 30352 9826 30359
rect 9876 30393 10646 30422
rect 9876 30359 9894 30393
rect 10062 30359 10152 30393
rect 10320 30359 10410 30393
rect 10578 30359 10646 30393
rect 8956 30342 9196 30352
rect 7506 30322 8296 30342
rect 7506 30321 8320 30322
rect 7504 30309 8324 30321
rect 7504 30249 7510 30309
rect 7544 30249 7768 30309
rect 7802 30249 8026 30309
rect 8060 30249 8284 30309
rect 8318 30249 8324 30309
rect 7504 30237 8324 30249
rect 8516 30247 8531 30322
rect 8586 30247 8606 30322
rect 8516 30237 8606 30247
rect 8746 30309 8886 30322
rect 8746 30249 8800 30309
rect 8834 30249 8886 30309
rect 6910 30202 7396 30212
rect 6910 30082 6966 30202
rect 7386 30082 7396 30202
rect 6910 30072 7396 30082
rect 7506 30152 8320 30237
rect 8746 30152 8886 30249
rect 9031 30309 9121 30342
rect 9876 30322 10646 30359
rect 9031 30249 9058 30309
rect 9092 30249 9121 30309
rect 9031 30232 9121 30249
rect 9266 30309 9406 30322
rect 9266 30249 9316 30309
rect 9350 30249 9406 30309
rect 9266 30152 9406 30249
rect 9551 30247 9561 30322
rect 9616 30247 9626 30322
rect 9551 30237 9626 30247
rect 9826 30309 10646 30322
rect 9826 30249 9832 30309
rect 9866 30249 10090 30309
rect 10124 30249 10348 30309
rect 10382 30249 10606 30309
rect 10640 30249 10646 30309
rect 9826 30152 10646 30249
rect 7506 30132 10646 30152
rect 7506 30062 7526 30132
rect 10626 30062 10646 30132
rect 7506 30042 10646 30062
rect 10836 29772 10946 31572
rect 6036 29752 10946 29772
rect 6036 29702 7466 29752
rect 10676 29702 10946 29752
rect 10986 29662 11036 31682
rect 5936 29592 7466 29662
rect 10676 29592 11036 29662
rect 5936 29572 11036 29592
rect 11136 29472 11216 31872
rect 5776 29372 11216 29472
rect 11256 29332 11336 32012
rect 12856 32012 13476 32092
rect 25848 32016 25948 32121
rect 26088 32297 26348 32316
rect 26088 32296 26141 32297
rect 26175 32296 26348 32297
rect 26088 32116 26108 32296
rect 26328 32116 26348 32296
rect 26088 32096 26348 32116
rect 26388 32296 27428 32316
rect 26388 32116 26408 32296
rect 26508 32116 27308 32296
rect 26388 32096 27308 32116
rect 26588 32076 27308 32096
rect 27388 32076 27428 32296
rect 26588 32056 27428 32076
rect 12856 31912 12956 32012
rect 13376 31912 13476 32012
rect 18368 31976 24068 31996
rect 13856 31912 14696 31952
rect 12716 31892 12976 31912
rect 11596 31732 11856 31752
rect 11596 31252 11616 31732
rect 11836 31252 11856 31732
rect 12716 31712 12736 31892
rect 12956 31712 12976 31892
rect 13356 31892 13616 31912
rect 12716 31701 12893 31712
rect 12927 31701 12976 31712
rect 12716 31692 12976 31701
rect 13145 31877 13191 31889
rect 13145 31701 13151 31877
rect 13185 31701 13191 31877
rect 12887 31689 12933 31692
rect 13145 31689 13191 31701
rect 13356 31712 13376 31892
rect 13596 31712 13616 31892
rect 13356 31701 13409 31712
rect 13443 31701 13616 31712
rect 13356 31692 13616 31701
rect 13656 31892 14396 31912
rect 13656 31712 13676 31892
rect 13776 31712 14396 31892
rect 13656 31692 14396 31712
rect 14476 31692 14696 31912
rect 13403 31689 13449 31692
rect 12943 31652 13135 31657
rect 13201 31652 13393 31657
rect 13856 31652 14696 31692
rect 18368 31936 20198 31976
rect 23408 31936 24068 31976
rect 12936 31651 13396 31652
rect 12936 31617 12955 31651
rect 13123 31617 13213 31651
rect 13381 31617 13396 31651
rect 12936 31552 13396 31617
rect 12936 31372 12956 31552
rect 13376 31372 13396 31552
rect 12936 31352 13396 31372
rect 11596 31232 11856 31252
rect 12936 31252 13396 31272
rect 12936 31072 12956 31252
rect 13376 31072 13396 31252
rect 12936 31006 13396 31072
rect 12936 30972 12955 31006
rect 13123 30972 13213 31006
rect 13381 30972 13396 31006
rect 12943 30966 13135 30972
rect 13201 30966 13393 30972
rect 13856 30932 14696 30972
rect 12716 30913 12976 30932
rect 12716 30912 12893 30913
rect 12927 30912 12976 30913
rect 12716 30732 12736 30912
rect 12956 30732 12976 30912
rect 12716 30712 12976 30732
rect 13116 30913 13216 30932
rect 13116 30737 13151 30913
rect 13185 30737 13216 30913
rect 13116 30632 13216 30737
rect 13356 30913 13616 30932
rect 13356 30912 13409 30913
rect 13443 30912 13616 30913
rect 13356 30732 13376 30912
rect 13596 30732 13616 30912
rect 13356 30712 13616 30732
rect 13656 30912 14696 30932
rect 13656 30732 13676 30912
rect 13776 30732 14576 30912
rect 13656 30712 14576 30732
rect 13856 30692 14576 30712
rect 14656 30692 14696 30912
rect 13856 30672 14696 30692
rect 12856 30552 13476 30632
rect 12856 30452 12956 30552
rect 13376 30452 13476 30552
rect 13856 30452 14696 30492
rect 12716 30432 12976 30452
rect 12716 30252 12736 30432
rect 12956 30252 12976 30432
rect 13356 30432 13616 30452
rect 12716 30241 12893 30252
rect 12927 30241 12976 30252
rect 12716 30232 12976 30241
rect 13145 30417 13191 30429
rect 13145 30241 13151 30417
rect 13185 30241 13191 30417
rect 12887 30229 12933 30232
rect 13145 30229 13191 30241
rect 13356 30252 13376 30432
rect 13596 30252 13616 30432
rect 13356 30241 13409 30252
rect 13443 30241 13616 30252
rect 13356 30232 13616 30241
rect 13656 30432 14396 30452
rect 13656 30252 13676 30432
rect 13776 30252 14396 30432
rect 13656 30232 14396 30252
rect 14476 30232 14696 30452
rect 13403 30229 13449 30232
rect 12943 30192 13135 30197
rect 13201 30192 13393 30197
rect 13856 30192 14696 30232
rect 12936 30191 13396 30192
rect 12936 30157 12955 30191
rect 13123 30157 13213 30191
rect 13381 30157 13396 30191
rect 11436 30132 11576 30152
rect 11436 29692 11456 30132
rect 11556 29692 11576 30132
rect 12936 30092 13396 30157
rect 12936 29912 12956 30092
rect 13376 29912 13396 30092
rect 12936 29892 13396 29912
rect 11436 29672 11576 29692
rect 12574 29552 13586 29572
rect 12574 29492 12596 29552
rect 13556 29541 13586 29552
rect 13557 29507 13586 29541
rect 13556 29492 13586 29507
rect 12574 29476 13586 29492
rect 5636 29272 11336 29332
rect 12216 29312 13216 29332
rect 11616 29273 11816 29292
rect 11616 29272 11658 29273
rect 11764 29272 11816 29273
rect 9536 29150 10696 29152
rect 9532 29132 10696 29150
rect 9532 29052 9556 29132
rect 10676 29052 10696 29132
rect 9532 29032 10696 29052
rect 9532 28980 10120 29032
rect 11616 29012 11636 29272
rect 9532 28874 9660 28980
rect 10057 28874 10120 28980
rect 9532 28838 10120 28874
rect 10836 28992 11636 29012
rect 10836 28812 10856 28992
rect 11796 28812 11816 29272
rect 12216 29132 12236 29312
rect 12416 29236 13216 29312
rect 12416 29202 12718 29236
rect 13206 29202 13216 29236
rect 12416 29132 13216 29202
rect 12216 29112 13216 29132
rect 13316 29312 13716 29332
rect 13316 29300 13516 29312
rect 13316 29136 13330 29300
rect 13378 29136 13516 29300
rect 13316 29132 13516 29136
rect 13696 29132 13716 29312
rect 18368 29256 18468 31936
rect 18508 31816 20198 31896
rect 23408 31816 23948 31896
rect 18508 31796 23948 31816
rect 18508 29396 18568 31796
rect 18668 31606 23768 31696
rect 18668 29586 18728 31606
rect 18768 31496 23678 31566
rect 18768 29696 18868 31496
rect 19642 31256 23378 31276
rect 19642 31236 20198 31256
rect 19642 31196 19748 31236
rect 19642 31176 20198 31196
rect 23358 31176 23378 31256
rect 19642 31156 23378 31176
rect 20238 31108 20298 31156
rect 20236 31096 20298 31108
rect 20488 31106 20548 31116
rect 20236 30920 20242 31096
rect 20276 30920 20298 31096
rect 20236 30908 20298 30920
rect 20448 31096 20598 31106
rect 20448 30986 20500 31096
rect 20534 30986 20598 31096
rect 20448 30926 20458 30986
rect 20568 30926 20598 30986
rect 20448 30920 20500 30926
rect 20534 30920 20598 30926
rect 20448 30916 20598 30920
rect 20708 31096 20838 31156
rect 21010 31106 21056 31108
rect 20708 30920 20758 31096
rect 20792 30920 20838 31096
rect 20708 30916 20838 30920
rect 20968 31096 21098 31106
rect 20968 30986 21016 31096
rect 21050 30986 21098 31096
rect 20968 30926 20978 30986
rect 21088 30926 21098 30986
rect 20968 30920 21016 30926
rect 21050 30920 21098 30926
rect 20968 30916 21098 30920
rect 21228 31096 21358 31156
rect 21228 30920 21274 31096
rect 21308 30920 21358 31096
rect 21228 30916 21358 30920
rect 21478 31096 21608 31116
rect 21478 30986 21532 31096
rect 21566 30986 21608 31096
rect 20238 30867 20298 30908
rect 20488 30906 20598 30916
rect 20752 30908 20798 30916
rect 21010 30908 21056 30916
rect 21268 30908 21314 30916
rect 20548 30867 20598 30906
rect 21478 30876 21488 30986
rect 21598 30876 21608 30986
rect 21738 31096 21868 31156
rect 22042 31106 22088 31108
rect 21738 30920 21790 31096
rect 21824 30920 21868 31096
rect 21738 30916 21868 30920
rect 21998 31096 22128 31106
rect 21998 30996 22048 31096
rect 22082 30996 22128 31096
rect 21998 30926 22008 30996
rect 22118 30926 22128 30996
rect 21998 30920 22048 30926
rect 22082 30920 22128 30926
rect 21998 30916 22128 30920
rect 22258 31096 22388 31156
rect 22258 30920 22306 31096
rect 22340 30920 22388 31096
rect 22258 30916 22388 30920
rect 22518 31096 22648 31116
rect 22518 30996 22564 31096
rect 22598 30996 22648 31096
rect 21784 30908 21830 30916
rect 22042 30908 22088 30916
rect 22300 30908 22346 30916
rect 21478 30867 21608 30876
rect 22518 30876 22528 30996
rect 22638 30876 22648 30996
rect 22778 31096 22908 31156
rect 23338 31108 23378 31156
rect 23074 31106 23120 31108
rect 22778 30920 22822 31096
rect 22856 30920 22908 31096
rect 22778 30916 22908 30920
rect 23028 31096 23158 31106
rect 23028 30996 23080 31096
rect 23114 30996 23158 31096
rect 23028 30926 23038 30996
rect 23148 30926 23158 30996
rect 23028 30920 23080 30926
rect 23114 30920 23158 30926
rect 23028 30916 23158 30920
rect 23332 31096 23378 31108
rect 23332 30920 23338 31096
rect 23372 30920 23378 31096
rect 22816 30908 22862 30916
rect 23074 30908 23120 30916
rect 23332 30908 23378 30920
rect 23338 30876 23378 30908
rect 22518 30867 22648 30876
rect 20238 30866 20484 30867
rect 20238 30861 20488 30866
rect 20548 30861 20742 30867
rect 20808 30861 21000 30867
rect 21066 30861 21258 30867
rect 21324 30861 21774 30867
rect 21840 30861 22032 30867
rect 22098 30861 22290 30867
rect 22356 30861 22806 30867
rect 22872 30861 23064 30867
rect 23128 30861 23378 30876
rect 20238 30827 20304 30861
rect 20472 30827 20488 30861
rect 20546 30827 20562 30861
rect 20730 30827 20820 30861
rect 20988 30827 21078 30861
rect 21246 30827 21336 30861
rect 21504 30827 21594 30861
rect 21762 30827 21852 30861
rect 22020 30827 22110 30861
rect 22278 30827 22368 30861
rect 22536 30827 22626 30861
rect 22794 30827 22884 30861
rect 23052 30827 23068 30861
rect 23128 30827 23142 30861
rect 23310 30827 23378 30861
rect 20238 30826 20488 30827
rect 20548 30826 20742 30827
rect 20292 30821 20484 30826
rect 20550 30821 20742 30826
rect 20808 30821 21000 30827
rect 21066 30821 21258 30827
rect 21324 30821 21516 30827
rect 21582 30821 21774 30827
rect 21840 30821 22032 30827
rect 22098 30821 22290 30827
rect 22356 30821 22548 30827
rect 22614 30821 22806 30827
rect 22872 30821 23064 30827
rect 23128 30826 23378 30827
rect 23130 30821 23322 30826
rect 20828 30776 20938 30786
rect 20550 30753 20742 30759
rect 20828 30753 20838 30776
rect 20546 30719 20562 30753
rect 20730 30719 20838 30753
rect 20550 30713 20742 30719
rect 20238 30681 20288 30686
rect 20236 30669 20288 30681
rect 20494 30676 20540 30681
rect 20236 30493 20242 30669
rect 20276 30493 20288 30669
rect 20236 30481 20288 30493
rect 20448 30669 20578 30676
rect 20448 30666 20500 30669
rect 20534 30666 20578 30669
rect 20448 30606 20458 30666
rect 20568 30606 20578 30666
rect 20448 30493 20500 30606
rect 20534 30493 20578 30606
rect 20752 30669 20798 30681
rect 20752 30576 20758 30669
rect 20448 30486 20578 30493
rect 20708 30556 20758 30576
rect 20792 30576 20798 30669
rect 20828 30616 20838 30719
rect 20928 30753 20938 30776
rect 22898 30776 22998 30786
rect 21324 30753 21516 30759
rect 21582 30753 21774 30759
rect 22356 30753 22548 30759
rect 22614 30753 22806 30759
rect 20928 30719 21336 30753
rect 21504 30719 21594 30753
rect 21762 30719 22368 30753
rect 22536 30719 22626 30753
rect 22794 30719 22810 30753
rect 20928 30616 20938 30719
rect 21324 30713 21516 30719
rect 21582 30713 21774 30719
rect 22356 30713 22548 30719
rect 22614 30713 22806 30719
rect 21010 30676 21056 30681
rect 21268 30676 21314 30681
rect 21526 30676 21572 30681
rect 21784 30676 21830 30681
rect 22042 30676 22088 30681
rect 22300 30676 22346 30681
rect 22558 30676 22604 30681
rect 20828 30606 20938 30616
rect 20968 30669 21098 30676
rect 20968 30666 21016 30669
rect 21050 30666 21098 30669
rect 20968 30606 20978 30666
rect 21088 30606 21098 30666
rect 20792 30556 20838 30576
rect 20708 30496 20718 30556
rect 20828 30496 20838 30556
rect 20708 30493 20758 30496
rect 20792 30493 20838 30496
rect 20708 30486 20838 30493
rect 20968 30493 21016 30606
rect 21050 30493 21098 30606
rect 20968 30486 21098 30493
rect 21228 30669 21358 30676
rect 21228 30556 21274 30669
rect 21308 30556 21358 30669
rect 21228 30496 21238 30556
rect 21348 30496 21358 30556
rect 21228 30493 21274 30496
rect 21308 30493 21358 30496
rect 21228 30486 21358 30493
rect 21478 30669 21608 30676
rect 21478 30666 21532 30669
rect 21566 30666 21608 30669
rect 21478 30606 21488 30666
rect 21598 30606 21608 30666
rect 21478 30493 21532 30606
rect 21566 30493 21608 30606
rect 21478 30486 21608 30493
rect 21748 30669 21878 30676
rect 21748 30556 21790 30669
rect 21824 30556 21878 30669
rect 21748 30496 21758 30556
rect 21868 30496 21878 30556
rect 21748 30493 21790 30496
rect 21824 30493 21878 30496
rect 21748 30486 21878 30493
rect 21998 30669 22128 30676
rect 21998 30666 22048 30669
rect 22082 30666 22128 30669
rect 21998 30606 22008 30666
rect 22118 30606 22128 30666
rect 21998 30493 22048 30606
rect 22082 30493 22128 30606
rect 21998 30486 22128 30493
rect 22258 30669 22388 30676
rect 22258 30556 22306 30669
rect 22340 30556 22388 30669
rect 22258 30496 22268 30556
rect 22378 30496 22388 30556
rect 22258 30493 22306 30496
rect 22340 30493 22388 30496
rect 22258 30486 22388 30493
rect 22518 30669 22648 30676
rect 22518 30666 22564 30669
rect 22598 30666 22648 30669
rect 22518 30606 22528 30666
rect 22638 30606 22648 30666
rect 22518 30493 22564 30606
rect 22598 30493 22648 30606
rect 22816 30669 22862 30681
rect 22816 30566 22822 30669
rect 22518 30486 22648 30493
rect 22768 30556 22822 30566
rect 22856 30566 22862 30669
rect 22898 30626 22908 30776
rect 22988 30626 22998 30776
rect 23074 30676 23120 30681
rect 22898 30596 22998 30626
rect 22856 30556 22898 30566
rect 22768 30496 22778 30556
rect 22888 30496 22898 30556
rect 22768 30493 22822 30496
rect 22856 30493 22898 30496
rect 22768 30486 22898 30493
rect 20494 30481 20540 30486
rect 20752 30481 20798 30486
rect 21010 30481 21056 30486
rect 21268 30481 21314 30486
rect 21526 30481 21572 30486
rect 21784 30481 21830 30486
rect 22042 30481 22088 30486
rect 22300 30481 22346 30486
rect 22558 30481 22604 30486
rect 22816 30481 22862 30486
rect 20238 30476 20288 30481
rect 20238 30449 20308 30476
rect 22928 30449 22998 30596
rect 23028 30669 23158 30676
rect 23028 30666 23080 30669
rect 23114 30666 23158 30669
rect 23028 30606 23038 30666
rect 23148 30606 23158 30666
rect 23028 30493 23080 30606
rect 23114 30493 23158 30606
rect 23028 30486 23158 30493
rect 23328 30669 23378 30686
rect 23328 30493 23338 30669
rect 23372 30493 23378 30669
rect 23074 30481 23120 30486
rect 23328 30476 23378 30493
rect 23298 30449 23378 30476
rect 20238 30446 20484 30449
rect 20238 30443 20488 30446
rect 20808 30443 21000 30449
rect 21066 30443 21258 30449
rect 21840 30443 22032 30449
rect 22098 30443 22290 30449
rect 22872 30443 23064 30449
rect 23130 30446 23378 30449
rect 23118 30443 23378 30446
rect 20238 30409 20304 30443
rect 20472 30409 20488 30443
rect 20804 30409 20820 30443
rect 20988 30409 21078 30443
rect 21246 30409 21852 30443
rect 22020 30409 22110 30443
rect 22278 30409 22884 30443
rect 23052 30409 23068 30443
rect 23118 30409 23142 30443
rect 23310 30409 23378 30443
rect 20238 30346 20488 30409
rect 20808 30403 21000 30409
rect 21066 30403 21258 30409
rect 21840 30403 22032 30409
rect 22098 30403 22290 30409
rect 22872 30403 23064 30409
rect 20238 30317 21008 30346
rect 21688 30336 21698 30366
rect 20238 30283 20304 30317
rect 20472 30283 20562 30317
rect 20730 30283 20820 30317
rect 20988 30283 21008 30317
rect 20238 30266 21008 30283
rect 21058 30317 21698 30336
rect 21918 30336 21928 30366
rect 23118 30346 23378 30409
rect 21918 30317 22558 30336
rect 21058 30283 21078 30317
rect 21246 30283 21336 30317
rect 21504 30283 21594 30317
rect 21762 30283 21852 30306
rect 22020 30283 22110 30317
rect 22278 30283 22368 30317
rect 22536 30283 22558 30317
rect 21058 30276 22558 30283
rect 22608 30317 23378 30346
rect 22608 30283 22626 30317
rect 22794 30283 22884 30317
rect 23052 30283 23142 30317
rect 23310 30283 23378 30317
rect 21688 30266 21928 30276
rect 20238 30246 21028 30266
rect 20238 30245 21052 30246
rect 20236 30233 21056 30245
rect 20236 30173 20242 30233
rect 20276 30173 20500 30233
rect 20534 30173 20758 30233
rect 20792 30173 21016 30233
rect 21050 30173 21056 30233
rect 20236 30161 21056 30173
rect 21248 30171 21263 30246
rect 21318 30171 21338 30246
rect 21248 30161 21338 30171
rect 21478 30233 21618 30246
rect 21478 30173 21532 30233
rect 21566 30173 21618 30233
rect 19642 30126 20128 30136
rect 19642 30006 19698 30126
rect 20118 30006 20128 30126
rect 19642 29996 20128 30006
rect 20238 30076 21052 30161
rect 21478 30076 21618 30173
rect 21763 30233 21853 30266
rect 22608 30246 23378 30283
rect 21763 30173 21790 30233
rect 21824 30173 21853 30233
rect 21763 30156 21853 30173
rect 21998 30233 22138 30246
rect 21998 30173 22048 30233
rect 22082 30173 22138 30233
rect 21998 30076 22138 30173
rect 22283 30171 22293 30246
rect 22348 30171 22358 30246
rect 22283 30161 22358 30171
rect 22558 30233 23378 30246
rect 22558 30173 22564 30233
rect 22598 30173 22822 30233
rect 22856 30173 23080 30233
rect 23114 30173 23338 30233
rect 23372 30173 23378 30233
rect 22558 30076 23378 30173
rect 20238 30056 23378 30076
rect 20238 29986 20258 30056
rect 23358 29986 23378 30056
rect 20238 29966 23378 29986
rect 23568 29696 23678 31496
rect 18768 29676 23678 29696
rect 18768 29626 20198 29676
rect 23408 29626 23678 29676
rect 23718 29586 23768 31606
rect 18668 29516 20198 29586
rect 23408 29516 23768 29586
rect 18668 29496 23768 29516
rect 23868 29396 23948 31796
rect 18508 29296 23948 29396
rect 23988 29256 24068 31936
rect 25588 31936 26208 32016
rect 25588 31836 25688 31936
rect 26108 31836 26208 31936
rect 26588 31836 27428 31876
rect 25448 31816 25708 31836
rect 24328 31656 24588 31676
rect 24328 31176 24348 31656
rect 24568 31176 24588 31656
rect 25448 31636 25468 31816
rect 25688 31636 25708 31816
rect 26088 31816 26348 31836
rect 25448 31625 25625 31636
rect 25659 31625 25708 31636
rect 25448 31616 25708 31625
rect 25877 31801 25923 31813
rect 25877 31625 25883 31801
rect 25917 31625 25923 31801
rect 25619 31613 25665 31616
rect 25877 31613 25923 31625
rect 26088 31636 26108 31816
rect 26328 31636 26348 31816
rect 26088 31625 26141 31636
rect 26175 31625 26348 31636
rect 26088 31616 26348 31625
rect 26388 31816 27128 31836
rect 26388 31636 26408 31816
rect 26508 31636 27128 31816
rect 26388 31616 27128 31636
rect 27208 31616 27428 31836
rect 26135 31613 26181 31616
rect 25675 31576 25867 31581
rect 25933 31576 26125 31581
rect 26588 31576 27428 31616
rect 25668 31575 26128 31576
rect 25668 31541 25687 31575
rect 25855 31541 25945 31575
rect 26113 31541 26128 31575
rect 25668 31476 26128 31541
rect 25668 31296 25688 31476
rect 26108 31296 26128 31476
rect 25668 31276 26128 31296
rect 24328 31156 24588 31176
rect 25668 31176 26128 31196
rect 25668 30996 25688 31176
rect 26108 30996 26128 31176
rect 25668 30930 26128 30996
rect 25668 30896 25687 30930
rect 25855 30896 25945 30930
rect 26113 30896 26128 30930
rect 25675 30890 25867 30896
rect 25933 30890 26125 30896
rect 26588 30856 27428 30896
rect 25448 30837 25708 30856
rect 25448 30836 25625 30837
rect 25659 30836 25708 30837
rect 25448 30656 25468 30836
rect 25688 30656 25708 30836
rect 25448 30636 25708 30656
rect 25848 30837 25948 30856
rect 25848 30661 25883 30837
rect 25917 30661 25948 30837
rect 25848 30556 25948 30661
rect 26088 30837 26348 30856
rect 26088 30836 26141 30837
rect 26175 30836 26348 30837
rect 26088 30656 26108 30836
rect 26328 30656 26348 30836
rect 26088 30636 26348 30656
rect 26388 30836 27428 30856
rect 26388 30656 26408 30836
rect 26508 30656 27308 30836
rect 26388 30636 27308 30656
rect 26588 30616 27308 30636
rect 27388 30616 27428 30836
rect 26588 30596 27428 30616
rect 25588 30476 26208 30556
rect 25588 30376 25688 30476
rect 26108 30376 26208 30476
rect 26588 30376 27428 30416
rect 25448 30356 25708 30376
rect 25448 30176 25468 30356
rect 25688 30176 25708 30356
rect 26088 30356 26348 30376
rect 25448 30165 25625 30176
rect 25659 30165 25708 30176
rect 25448 30156 25708 30165
rect 25877 30341 25923 30353
rect 25877 30165 25883 30341
rect 25917 30165 25923 30341
rect 25619 30153 25665 30156
rect 25877 30153 25923 30165
rect 26088 30176 26108 30356
rect 26328 30176 26348 30356
rect 26088 30165 26141 30176
rect 26175 30165 26348 30176
rect 26088 30156 26348 30165
rect 26388 30356 27128 30376
rect 26388 30176 26408 30356
rect 26508 30176 27128 30356
rect 26388 30156 27128 30176
rect 27208 30156 27428 30376
rect 26135 30153 26181 30156
rect 25675 30116 25867 30121
rect 25933 30116 26125 30121
rect 26588 30116 27428 30156
rect 25668 30115 26128 30116
rect 25668 30081 25687 30115
rect 25855 30081 25945 30115
rect 26113 30081 26128 30115
rect 24168 30056 24308 30076
rect 24168 29616 24188 30056
rect 24288 29616 24308 30056
rect 25668 30016 26128 30081
rect 25668 29836 25688 30016
rect 26108 29836 26128 30016
rect 25668 29816 26128 29836
rect 24168 29596 24308 29616
rect 25306 29476 26318 29496
rect 25306 29416 25328 29476
rect 26288 29465 26318 29476
rect 26289 29431 26318 29465
rect 26288 29416 26318 29431
rect 25306 29400 26318 29416
rect 18368 29196 24068 29256
rect 24948 29236 25948 29256
rect 24348 29197 24548 29216
rect 24348 29196 24390 29197
rect 24496 29196 24548 29197
rect 13316 29112 13716 29132
rect 22268 29074 23428 29076
rect 22264 29056 23428 29074
rect 12574 29012 13586 29028
rect 12574 28952 12596 29012
rect 13576 28952 13586 29012
rect 12574 28932 13586 28952
rect 22264 28976 22288 29056
rect 23408 28976 23428 29056
rect 22264 28956 23428 28976
rect 10836 28792 11816 28812
rect 22264 28904 22852 28956
rect 24348 28936 24368 29196
rect 22264 28798 22392 28904
rect 22789 28798 22852 28904
rect 22264 28762 22852 28798
rect 23568 28916 24368 28936
rect 23568 28736 23588 28916
rect 24528 28736 24548 29196
rect 24948 29056 24968 29236
rect 25148 29160 25948 29236
rect 25148 29126 25450 29160
rect 25938 29126 25948 29160
rect 25148 29056 25948 29126
rect 24948 29036 25948 29056
rect 26048 29236 26448 29256
rect 26048 29224 26248 29236
rect 26048 29060 26062 29224
rect 26110 29060 26248 29224
rect 26048 29056 26248 29060
rect 26428 29056 26448 29236
rect 26048 29036 26448 29056
rect 25306 28936 26318 28952
rect 25306 28876 25328 28936
rect 26308 28876 26318 28936
rect 25306 28856 26318 28876
rect 23568 28716 24548 28736
rect 13056 26008 13516 26028
rect 13056 25828 13076 26008
rect 13496 25828 13516 26008
rect 13056 25762 13516 25828
rect 13056 25728 13075 25762
rect 13243 25728 13333 25762
rect 13501 25728 13516 25762
rect 25764 25878 26224 25898
rect 13063 25722 13255 25728
rect 13321 25722 13513 25728
rect 13976 25688 14816 25728
rect 12836 25669 13096 25688
rect 12836 25668 13013 25669
rect 13047 25668 13096 25669
rect 12836 25488 12856 25668
rect 13076 25488 13096 25668
rect 12836 25468 13096 25488
rect 13236 25669 13336 25688
rect 13236 25493 13271 25669
rect 13305 25493 13336 25669
rect 13236 25388 13336 25493
rect 13476 25669 13736 25688
rect 13476 25668 13529 25669
rect 13563 25668 13736 25669
rect 13476 25488 13496 25668
rect 13716 25488 13736 25668
rect 13476 25468 13736 25488
rect 13776 25668 14816 25688
rect 13776 25488 13796 25668
rect 13896 25488 14696 25668
rect 13776 25468 14696 25488
rect 13976 25448 14696 25468
rect 14776 25448 14816 25668
rect 25764 25698 25784 25878
rect 26204 25698 26224 25878
rect 25764 25632 26224 25698
rect 25764 25598 25783 25632
rect 25951 25598 26041 25632
rect 26209 25598 26224 25632
rect 25771 25592 25963 25598
rect 26029 25592 26221 25598
rect 26684 25558 27524 25598
rect 13976 25428 14816 25448
rect 25544 25539 25804 25558
rect 25544 25538 25721 25539
rect 25755 25538 25804 25539
rect 5756 25348 11456 25368
rect 5756 25308 7586 25348
rect 10796 25308 11456 25348
rect 5756 22628 5856 25308
rect 5896 25188 7586 25268
rect 10796 25188 11336 25268
rect 5896 25168 11336 25188
rect 5896 22768 5956 25168
rect 6056 24978 11156 25068
rect 6056 22958 6116 24978
rect 6156 24868 11066 24938
rect 6156 23068 6256 24868
rect 7030 24628 10766 24648
rect 7030 24608 7586 24628
rect 7030 24568 7136 24608
rect 7030 24548 7586 24568
rect 10746 24548 10766 24628
rect 7030 24528 10766 24548
rect 7626 24480 7686 24528
rect 7624 24468 7686 24480
rect 7876 24478 7936 24488
rect 7624 24292 7630 24468
rect 7664 24292 7686 24468
rect 7624 24280 7686 24292
rect 7836 24468 7986 24478
rect 7836 24358 7888 24468
rect 7922 24358 7986 24468
rect 7836 24298 7846 24358
rect 7956 24298 7986 24358
rect 7836 24292 7888 24298
rect 7922 24292 7986 24298
rect 7836 24288 7986 24292
rect 8096 24468 8226 24528
rect 8398 24478 8444 24480
rect 8096 24292 8146 24468
rect 8180 24292 8226 24468
rect 8096 24288 8226 24292
rect 8356 24468 8486 24478
rect 8356 24358 8404 24468
rect 8438 24358 8486 24468
rect 8356 24298 8366 24358
rect 8476 24298 8486 24358
rect 8356 24292 8404 24298
rect 8438 24292 8486 24298
rect 8356 24288 8486 24292
rect 8616 24468 8746 24528
rect 8616 24292 8662 24468
rect 8696 24292 8746 24468
rect 8616 24288 8746 24292
rect 8866 24468 8996 24488
rect 8866 24358 8920 24468
rect 8954 24358 8996 24468
rect 7626 24239 7686 24280
rect 7876 24278 7986 24288
rect 8140 24280 8186 24288
rect 8398 24280 8444 24288
rect 8656 24280 8702 24288
rect 7936 24239 7986 24278
rect 8866 24248 8876 24358
rect 8986 24248 8996 24358
rect 9126 24468 9256 24528
rect 9430 24478 9476 24480
rect 9126 24292 9178 24468
rect 9212 24292 9256 24468
rect 9126 24288 9256 24292
rect 9386 24468 9516 24478
rect 9386 24368 9436 24468
rect 9470 24368 9516 24468
rect 9386 24298 9396 24368
rect 9506 24298 9516 24368
rect 9386 24292 9436 24298
rect 9470 24292 9516 24298
rect 9386 24288 9516 24292
rect 9646 24468 9776 24528
rect 9646 24292 9694 24468
rect 9728 24292 9776 24468
rect 9646 24288 9776 24292
rect 9906 24468 10036 24488
rect 9906 24368 9952 24468
rect 9986 24368 10036 24468
rect 9172 24280 9218 24288
rect 9430 24280 9476 24288
rect 9688 24280 9734 24288
rect 8866 24239 8996 24248
rect 9906 24248 9916 24368
rect 10026 24248 10036 24368
rect 10166 24468 10296 24528
rect 10726 24480 10766 24528
rect 10462 24478 10508 24480
rect 10166 24292 10210 24468
rect 10244 24292 10296 24468
rect 10166 24288 10296 24292
rect 10416 24468 10546 24478
rect 10416 24368 10468 24468
rect 10502 24368 10546 24468
rect 10416 24298 10426 24368
rect 10536 24298 10546 24368
rect 10416 24292 10468 24298
rect 10502 24292 10546 24298
rect 10416 24288 10546 24292
rect 10720 24468 10766 24480
rect 10720 24292 10726 24468
rect 10760 24292 10766 24468
rect 10204 24280 10250 24288
rect 10462 24280 10508 24288
rect 10720 24280 10766 24292
rect 10726 24248 10766 24280
rect 9906 24239 10036 24248
rect 7626 24238 7872 24239
rect 7626 24233 7876 24238
rect 7936 24233 8130 24239
rect 8196 24233 8388 24239
rect 8454 24233 8646 24239
rect 8712 24233 9162 24239
rect 9228 24233 9420 24239
rect 9486 24233 9678 24239
rect 9744 24233 10194 24239
rect 10260 24233 10452 24239
rect 10516 24233 10766 24248
rect 7626 24199 7692 24233
rect 7860 24199 7876 24233
rect 7934 24199 7950 24233
rect 8118 24199 8208 24233
rect 8376 24199 8466 24233
rect 8634 24199 8724 24233
rect 8892 24199 8982 24233
rect 9150 24199 9240 24233
rect 9408 24199 9498 24233
rect 9666 24199 9756 24233
rect 9924 24199 10014 24233
rect 10182 24199 10272 24233
rect 10440 24199 10456 24233
rect 10516 24199 10530 24233
rect 10698 24199 10766 24233
rect 7626 24198 7876 24199
rect 7936 24198 8130 24199
rect 7680 24193 7872 24198
rect 7938 24193 8130 24198
rect 8196 24193 8388 24199
rect 8454 24193 8646 24199
rect 8712 24193 8904 24199
rect 8970 24193 9162 24199
rect 9228 24193 9420 24199
rect 9486 24193 9678 24199
rect 9744 24193 9936 24199
rect 10002 24193 10194 24199
rect 10260 24193 10452 24199
rect 10516 24198 10766 24199
rect 10518 24193 10710 24198
rect 8216 24148 8326 24158
rect 7938 24125 8130 24131
rect 8216 24125 8226 24148
rect 7934 24091 7950 24125
rect 8118 24091 8226 24125
rect 7938 24085 8130 24091
rect 7626 24053 7676 24058
rect 7624 24041 7676 24053
rect 7882 24048 7928 24053
rect 7624 23865 7630 24041
rect 7664 23865 7676 24041
rect 7624 23853 7676 23865
rect 7836 24041 7966 24048
rect 7836 24038 7888 24041
rect 7922 24038 7966 24041
rect 7836 23978 7846 24038
rect 7956 23978 7966 24038
rect 7836 23865 7888 23978
rect 7922 23865 7966 23978
rect 8140 24041 8186 24053
rect 8140 23948 8146 24041
rect 7836 23858 7966 23865
rect 8096 23928 8146 23948
rect 8180 23948 8186 24041
rect 8216 23988 8226 24091
rect 8316 24125 8326 24148
rect 10286 24148 10386 24158
rect 8712 24125 8904 24131
rect 8970 24125 9162 24131
rect 9744 24125 9936 24131
rect 10002 24125 10194 24131
rect 8316 24091 8724 24125
rect 8892 24091 8982 24125
rect 9150 24091 9756 24125
rect 9924 24091 10014 24125
rect 10182 24091 10198 24125
rect 8316 23988 8326 24091
rect 8712 24085 8904 24091
rect 8970 24085 9162 24091
rect 9744 24085 9936 24091
rect 10002 24085 10194 24091
rect 8398 24048 8444 24053
rect 8656 24048 8702 24053
rect 8914 24048 8960 24053
rect 9172 24048 9218 24053
rect 9430 24048 9476 24053
rect 9688 24048 9734 24053
rect 9946 24048 9992 24053
rect 8216 23978 8326 23988
rect 8356 24041 8486 24048
rect 8356 24038 8404 24041
rect 8438 24038 8486 24041
rect 8356 23978 8366 24038
rect 8476 23978 8486 24038
rect 8180 23928 8226 23948
rect 8096 23868 8106 23928
rect 8216 23868 8226 23928
rect 8096 23865 8146 23868
rect 8180 23865 8226 23868
rect 8096 23858 8226 23865
rect 8356 23865 8404 23978
rect 8438 23865 8486 23978
rect 8356 23858 8486 23865
rect 8616 24041 8746 24048
rect 8616 23928 8662 24041
rect 8696 23928 8746 24041
rect 8616 23868 8626 23928
rect 8736 23868 8746 23928
rect 8616 23865 8662 23868
rect 8696 23865 8746 23868
rect 8616 23858 8746 23865
rect 8866 24041 8996 24048
rect 8866 24038 8920 24041
rect 8954 24038 8996 24041
rect 8866 23978 8876 24038
rect 8986 23978 8996 24038
rect 8866 23865 8920 23978
rect 8954 23865 8996 23978
rect 8866 23858 8996 23865
rect 9136 24041 9266 24048
rect 9136 23928 9178 24041
rect 9212 23928 9266 24041
rect 9136 23868 9146 23928
rect 9256 23868 9266 23928
rect 9136 23865 9178 23868
rect 9212 23865 9266 23868
rect 9136 23858 9266 23865
rect 9386 24041 9516 24048
rect 9386 24038 9436 24041
rect 9470 24038 9516 24041
rect 9386 23978 9396 24038
rect 9506 23978 9516 24038
rect 9386 23865 9436 23978
rect 9470 23865 9516 23978
rect 9386 23858 9516 23865
rect 9646 24041 9776 24048
rect 9646 23928 9694 24041
rect 9728 23928 9776 24041
rect 9646 23868 9656 23928
rect 9766 23868 9776 23928
rect 9646 23865 9694 23868
rect 9728 23865 9776 23868
rect 9646 23858 9776 23865
rect 9906 24041 10036 24048
rect 9906 24038 9952 24041
rect 9986 24038 10036 24041
rect 9906 23978 9916 24038
rect 10026 23978 10036 24038
rect 9906 23865 9952 23978
rect 9986 23865 10036 23978
rect 10204 24041 10250 24053
rect 10204 23938 10210 24041
rect 9906 23858 10036 23865
rect 10156 23928 10210 23938
rect 10244 23938 10250 24041
rect 10286 23998 10296 24148
rect 10376 23998 10386 24148
rect 10462 24048 10508 24053
rect 10286 23968 10386 23998
rect 10244 23928 10286 23938
rect 10156 23868 10166 23928
rect 10276 23868 10286 23928
rect 10156 23865 10210 23868
rect 10244 23865 10286 23868
rect 10156 23858 10286 23865
rect 7882 23853 7928 23858
rect 8140 23853 8186 23858
rect 8398 23853 8444 23858
rect 8656 23853 8702 23858
rect 8914 23853 8960 23858
rect 9172 23853 9218 23858
rect 9430 23853 9476 23858
rect 9688 23853 9734 23858
rect 9946 23853 9992 23858
rect 10204 23853 10250 23858
rect 7626 23848 7676 23853
rect 7626 23821 7696 23848
rect 10316 23821 10386 23968
rect 10416 24041 10546 24048
rect 10416 24038 10468 24041
rect 10502 24038 10546 24041
rect 10416 23978 10426 24038
rect 10536 23978 10546 24038
rect 10416 23865 10468 23978
rect 10502 23865 10546 23978
rect 10416 23858 10546 23865
rect 10716 24041 10766 24058
rect 10716 23865 10726 24041
rect 10760 23865 10766 24041
rect 10462 23853 10508 23858
rect 10716 23848 10766 23865
rect 10686 23821 10766 23848
rect 7626 23818 7872 23821
rect 7626 23815 7876 23818
rect 8196 23815 8388 23821
rect 8454 23815 8646 23821
rect 9228 23815 9420 23821
rect 9486 23815 9678 23821
rect 10260 23815 10452 23821
rect 10518 23818 10766 23821
rect 10506 23815 10766 23818
rect 7626 23781 7692 23815
rect 7860 23781 7876 23815
rect 8192 23781 8208 23815
rect 8376 23781 8466 23815
rect 8634 23781 9240 23815
rect 9408 23781 9498 23815
rect 9666 23781 10272 23815
rect 10440 23781 10456 23815
rect 10506 23781 10530 23815
rect 10698 23781 10766 23815
rect 7626 23718 7876 23781
rect 8196 23775 8388 23781
rect 8454 23775 8646 23781
rect 9228 23775 9420 23781
rect 9486 23775 9678 23781
rect 10260 23775 10452 23781
rect 7626 23689 8396 23718
rect 9076 23708 9086 23738
rect 7626 23655 7692 23689
rect 7860 23655 7950 23689
rect 8118 23655 8208 23689
rect 8376 23655 8396 23689
rect 7626 23638 8396 23655
rect 8446 23689 9086 23708
rect 9306 23708 9316 23738
rect 10506 23718 10766 23781
rect 9306 23689 9946 23708
rect 8446 23655 8466 23689
rect 8634 23655 8724 23689
rect 8892 23655 8982 23689
rect 9150 23655 9240 23678
rect 9408 23655 9498 23689
rect 9666 23655 9756 23689
rect 9924 23655 9946 23689
rect 8446 23648 9946 23655
rect 9996 23689 10766 23718
rect 9996 23655 10014 23689
rect 10182 23655 10272 23689
rect 10440 23655 10530 23689
rect 10698 23655 10766 23689
rect 9076 23638 9316 23648
rect 7626 23618 8416 23638
rect 7626 23617 8440 23618
rect 7624 23605 8444 23617
rect 7624 23545 7630 23605
rect 7664 23545 7888 23605
rect 7922 23545 8146 23605
rect 8180 23545 8404 23605
rect 8438 23545 8444 23605
rect 7624 23533 8444 23545
rect 8636 23543 8651 23618
rect 8706 23543 8726 23618
rect 8636 23533 8726 23543
rect 8866 23605 9006 23618
rect 8866 23545 8920 23605
rect 8954 23545 9006 23605
rect 7030 23498 7516 23508
rect 7030 23378 7086 23498
rect 7506 23378 7516 23498
rect 7030 23368 7516 23378
rect 7626 23448 8440 23533
rect 8866 23448 9006 23545
rect 9151 23605 9241 23638
rect 9996 23618 10766 23655
rect 9151 23545 9178 23605
rect 9212 23545 9241 23605
rect 9151 23528 9241 23545
rect 9386 23605 9526 23618
rect 9386 23545 9436 23605
rect 9470 23545 9526 23605
rect 9386 23448 9526 23545
rect 9671 23543 9681 23618
rect 9736 23543 9746 23618
rect 9671 23533 9746 23543
rect 9946 23605 10766 23618
rect 9946 23545 9952 23605
rect 9986 23545 10210 23605
rect 10244 23545 10468 23605
rect 10502 23545 10726 23605
rect 10760 23545 10766 23605
rect 9946 23448 10766 23545
rect 7626 23428 10766 23448
rect 7626 23358 7646 23428
rect 10746 23358 10766 23428
rect 7626 23338 10766 23358
rect 10956 23068 11066 24868
rect 6156 23048 11066 23068
rect 6156 22998 7586 23048
rect 10796 22998 11066 23048
rect 11106 22958 11156 24978
rect 6056 22888 7586 22958
rect 10796 22888 11156 22958
rect 6056 22868 11156 22888
rect 11256 22768 11336 25168
rect 5896 22668 11336 22768
rect 11376 22628 11456 25308
rect 12976 25308 13596 25388
rect 25544 25358 25564 25538
rect 25784 25358 25804 25538
rect 25544 25338 25804 25358
rect 25944 25539 26044 25558
rect 25944 25363 25979 25539
rect 26013 25363 26044 25539
rect 12976 25208 13076 25308
rect 13496 25208 13596 25308
rect 25944 25258 26044 25363
rect 26184 25539 26444 25558
rect 26184 25538 26237 25539
rect 26271 25538 26444 25539
rect 26184 25358 26204 25538
rect 26424 25358 26444 25538
rect 26184 25338 26444 25358
rect 26484 25538 27524 25558
rect 26484 25358 26504 25538
rect 26604 25358 27404 25538
rect 26484 25338 27404 25358
rect 26684 25318 27404 25338
rect 27484 25318 27524 25538
rect 26684 25298 27524 25318
rect 13976 25208 14816 25248
rect 12836 25188 13096 25208
rect 11716 25028 11976 25048
rect 11716 24548 11736 25028
rect 11956 24548 11976 25028
rect 12836 25008 12856 25188
rect 13076 25008 13096 25188
rect 13476 25188 13736 25208
rect 12836 24997 13013 25008
rect 13047 24997 13096 25008
rect 12836 24988 13096 24997
rect 13265 25173 13311 25185
rect 13265 24997 13271 25173
rect 13305 24997 13311 25173
rect 13007 24985 13053 24988
rect 13265 24985 13311 24997
rect 13476 25008 13496 25188
rect 13716 25008 13736 25188
rect 13476 24997 13529 25008
rect 13563 24997 13736 25008
rect 13476 24988 13736 24997
rect 13776 25188 14516 25208
rect 13776 25008 13796 25188
rect 13896 25008 14516 25188
rect 13776 24988 14516 25008
rect 14596 24988 14816 25208
rect 13523 24985 13569 24988
rect 13063 24948 13255 24953
rect 13321 24948 13513 24953
rect 13976 24948 14816 24988
rect 18464 25218 24164 25238
rect 18464 25178 20294 25218
rect 23504 25178 24164 25218
rect 13056 24947 13516 24948
rect 13056 24913 13075 24947
rect 13243 24913 13333 24947
rect 13501 24913 13516 24947
rect 13056 24848 13516 24913
rect 13056 24668 13076 24848
rect 13496 24668 13516 24848
rect 13056 24648 13516 24668
rect 11716 24528 11976 24548
rect 13056 24548 13516 24568
rect 13056 24368 13076 24548
rect 13496 24368 13516 24548
rect 13056 24302 13516 24368
rect 13056 24268 13075 24302
rect 13243 24268 13333 24302
rect 13501 24268 13516 24302
rect 13063 24262 13255 24268
rect 13321 24262 13513 24268
rect 13976 24228 14816 24268
rect 12836 24209 13096 24228
rect 12836 24208 13013 24209
rect 13047 24208 13096 24209
rect 12836 24028 12856 24208
rect 13076 24028 13096 24208
rect 12836 24008 13096 24028
rect 13236 24209 13336 24228
rect 13236 24033 13271 24209
rect 13305 24033 13336 24209
rect 13236 23928 13336 24033
rect 13476 24209 13736 24228
rect 13476 24208 13529 24209
rect 13563 24208 13736 24209
rect 13476 24028 13496 24208
rect 13716 24028 13736 24208
rect 13476 24008 13736 24028
rect 13776 24208 14816 24228
rect 13776 24028 13796 24208
rect 13896 24028 14696 24208
rect 13776 24008 14696 24028
rect 13976 23988 14696 24008
rect 14776 23988 14816 24208
rect 13976 23968 14816 23988
rect 12976 23848 13596 23928
rect 12976 23748 13076 23848
rect 13496 23748 13596 23848
rect 13976 23748 14816 23788
rect 12836 23728 13096 23748
rect 12836 23548 12856 23728
rect 13076 23548 13096 23728
rect 13476 23728 13736 23748
rect 12836 23537 13013 23548
rect 13047 23537 13096 23548
rect 12836 23528 13096 23537
rect 13265 23713 13311 23725
rect 13265 23537 13271 23713
rect 13305 23537 13311 23713
rect 13007 23525 13053 23528
rect 13265 23525 13311 23537
rect 13476 23548 13496 23728
rect 13716 23548 13736 23728
rect 13476 23537 13529 23548
rect 13563 23537 13736 23548
rect 13476 23528 13736 23537
rect 13776 23728 14516 23748
rect 13776 23548 13796 23728
rect 13896 23548 14516 23728
rect 13776 23528 14516 23548
rect 14596 23528 14816 23748
rect 13523 23525 13569 23528
rect 13063 23488 13255 23493
rect 13321 23488 13513 23493
rect 13976 23488 14816 23528
rect 13056 23487 13516 23488
rect 13056 23453 13075 23487
rect 13243 23453 13333 23487
rect 13501 23453 13516 23487
rect 11556 23428 11696 23448
rect 11556 22988 11576 23428
rect 11676 22988 11696 23428
rect 13056 23388 13516 23453
rect 13056 23208 13076 23388
rect 13496 23208 13516 23388
rect 13056 23188 13516 23208
rect 11556 22968 11696 22988
rect 12694 22848 13706 22868
rect 12694 22788 12716 22848
rect 13676 22837 13706 22848
rect 13677 22803 13706 22837
rect 13676 22788 13706 22803
rect 12694 22772 13706 22788
rect 5756 22568 11456 22628
rect 12336 22608 13336 22628
rect 11736 22569 11936 22588
rect 11736 22568 11778 22569
rect 11884 22568 11936 22569
rect 9656 22446 10816 22448
rect 9652 22428 10816 22446
rect 9652 22348 9676 22428
rect 10796 22348 10816 22428
rect 9652 22328 10816 22348
rect 9652 22276 10240 22328
rect 11736 22308 11756 22568
rect 9652 22170 9780 22276
rect 10177 22170 10240 22276
rect 9652 22134 10240 22170
rect 10956 22288 11756 22308
rect 10956 22108 10976 22288
rect 11916 22108 11936 22568
rect 12336 22428 12356 22608
rect 12536 22532 13336 22608
rect 12536 22498 12838 22532
rect 13326 22498 13336 22532
rect 12536 22428 13336 22498
rect 12336 22408 13336 22428
rect 13436 22608 13836 22628
rect 13436 22596 13636 22608
rect 13436 22432 13450 22596
rect 13498 22432 13636 22596
rect 13436 22428 13636 22432
rect 13816 22428 13836 22608
rect 18464 22498 18564 25178
rect 18604 25058 20294 25138
rect 23504 25058 24044 25138
rect 18604 25038 24044 25058
rect 18604 22638 18664 25038
rect 18764 24848 23864 24938
rect 18764 22828 18824 24848
rect 18864 24738 23774 24808
rect 18864 22938 18964 24738
rect 19738 24498 23474 24518
rect 19738 24478 20294 24498
rect 19738 24438 19844 24478
rect 19738 24418 20294 24438
rect 23454 24418 23474 24498
rect 19738 24398 23474 24418
rect 20334 24350 20394 24398
rect 20332 24338 20394 24350
rect 20584 24348 20644 24358
rect 20332 24162 20338 24338
rect 20372 24162 20394 24338
rect 20332 24150 20394 24162
rect 20544 24338 20694 24348
rect 20544 24228 20596 24338
rect 20630 24228 20694 24338
rect 20544 24168 20554 24228
rect 20664 24168 20694 24228
rect 20544 24162 20596 24168
rect 20630 24162 20694 24168
rect 20544 24158 20694 24162
rect 20804 24338 20934 24398
rect 21106 24348 21152 24350
rect 20804 24162 20854 24338
rect 20888 24162 20934 24338
rect 20804 24158 20934 24162
rect 21064 24338 21194 24348
rect 21064 24228 21112 24338
rect 21146 24228 21194 24338
rect 21064 24168 21074 24228
rect 21184 24168 21194 24228
rect 21064 24162 21112 24168
rect 21146 24162 21194 24168
rect 21064 24158 21194 24162
rect 21324 24338 21454 24398
rect 21324 24162 21370 24338
rect 21404 24162 21454 24338
rect 21324 24158 21454 24162
rect 21574 24338 21704 24358
rect 21574 24228 21628 24338
rect 21662 24228 21704 24338
rect 20334 24109 20394 24150
rect 20584 24148 20694 24158
rect 20848 24150 20894 24158
rect 21106 24150 21152 24158
rect 21364 24150 21410 24158
rect 20644 24109 20694 24148
rect 21574 24118 21584 24228
rect 21694 24118 21704 24228
rect 21834 24338 21964 24398
rect 22138 24348 22184 24350
rect 21834 24162 21886 24338
rect 21920 24162 21964 24338
rect 21834 24158 21964 24162
rect 22094 24338 22224 24348
rect 22094 24238 22144 24338
rect 22178 24238 22224 24338
rect 22094 24168 22104 24238
rect 22214 24168 22224 24238
rect 22094 24162 22144 24168
rect 22178 24162 22224 24168
rect 22094 24158 22224 24162
rect 22354 24338 22484 24398
rect 22354 24162 22402 24338
rect 22436 24162 22484 24338
rect 22354 24158 22484 24162
rect 22614 24338 22744 24358
rect 22614 24238 22660 24338
rect 22694 24238 22744 24338
rect 21880 24150 21926 24158
rect 22138 24150 22184 24158
rect 22396 24150 22442 24158
rect 21574 24109 21704 24118
rect 22614 24118 22624 24238
rect 22734 24118 22744 24238
rect 22874 24338 23004 24398
rect 23434 24350 23474 24398
rect 23170 24348 23216 24350
rect 22874 24162 22918 24338
rect 22952 24162 23004 24338
rect 22874 24158 23004 24162
rect 23124 24338 23254 24348
rect 23124 24238 23176 24338
rect 23210 24238 23254 24338
rect 23124 24168 23134 24238
rect 23244 24168 23254 24238
rect 23124 24162 23176 24168
rect 23210 24162 23254 24168
rect 23124 24158 23254 24162
rect 23428 24338 23474 24350
rect 23428 24162 23434 24338
rect 23468 24162 23474 24338
rect 22912 24150 22958 24158
rect 23170 24150 23216 24158
rect 23428 24150 23474 24162
rect 23434 24118 23474 24150
rect 22614 24109 22744 24118
rect 20334 24108 20580 24109
rect 20334 24103 20584 24108
rect 20644 24103 20838 24109
rect 20904 24103 21096 24109
rect 21162 24103 21354 24109
rect 21420 24103 21870 24109
rect 21936 24103 22128 24109
rect 22194 24103 22386 24109
rect 22452 24103 22902 24109
rect 22968 24103 23160 24109
rect 23224 24103 23474 24118
rect 20334 24069 20400 24103
rect 20568 24069 20584 24103
rect 20642 24069 20658 24103
rect 20826 24069 20916 24103
rect 21084 24069 21174 24103
rect 21342 24069 21432 24103
rect 21600 24069 21690 24103
rect 21858 24069 21948 24103
rect 22116 24069 22206 24103
rect 22374 24069 22464 24103
rect 22632 24069 22722 24103
rect 22890 24069 22980 24103
rect 23148 24069 23164 24103
rect 23224 24069 23238 24103
rect 23406 24069 23474 24103
rect 20334 24068 20584 24069
rect 20644 24068 20838 24069
rect 20388 24063 20580 24068
rect 20646 24063 20838 24068
rect 20904 24063 21096 24069
rect 21162 24063 21354 24069
rect 21420 24063 21612 24069
rect 21678 24063 21870 24069
rect 21936 24063 22128 24069
rect 22194 24063 22386 24069
rect 22452 24063 22644 24069
rect 22710 24063 22902 24069
rect 22968 24063 23160 24069
rect 23224 24068 23474 24069
rect 23226 24063 23418 24068
rect 20924 24018 21034 24028
rect 20646 23995 20838 24001
rect 20924 23995 20934 24018
rect 20642 23961 20658 23995
rect 20826 23961 20934 23995
rect 20646 23955 20838 23961
rect 20334 23923 20384 23928
rect 20332 23911 20384 23923
rect 20590 23918 20636 23923
rect 20332 23735 20338 23911
rect 20372 23735 20384 23911
rect 20332 23723 20384 23735
rect 20544 23911 20674 23918
rect 20544 23908 20596 23911
rect 20630 23908 20674 23911
rect 20544 23848 20554 23908
rect 20664 23848 20674 23908
rect 20544 23735 20596 23848
rect 20630 23735 20674 23848
rect 20848 23911 20894 23923
rect 20848 23818 20854 23911
rect 20544 23728 20674 23735
rect 20804 23798 20854 23818
rect 20888 23818 20894 23911
rect 20924 23858 20934 23961
rect 21024 23995 21034 24018
rect 22994 24018 23094 24028
rect 21420 23995 21612 24001
rect 21678 23995 21870 24001
rect 22452 23995 22644 24001
rect 22710 23995 22902 24001
rect 21024 23961 21432 23995
rect 21600 23961 21690 23995
rect 21858 23961 22464 23995
rect 22632 23961 22722 23995
rect 22890 23961 22906 23995
rect 21024 23858 21034 23961
rect 21420 23955 21612 23961
rect 21678 23955 21870 23961
rect 22452 23955 22644 23961
rect 22710 23955 22902 23961
rect 21106 23918 21152 23923
rect 21364 23918 21410 23923
rect 21622 23918 21668 23923
rect 21880 23918 21926 23923
rect 22138 23918 22184 23923
rect 22396 23918 22442 23923
rect 22654 23918 22700 23923
rect 20924 23848 21034 23858
rect 21064 23911 21194 23918
rect 21064 23908 21112 23911
rect 21146 23908 21194 23911
rect 21064 23848 21074 23908
rect 21184 23848 21194 23908
rect 20888 23798 20934 23818
rect 20804 23738 20814 23798
rect 20924 23738 20934 23798
rect 20804 23735 20854 23738
rect 20888 23735 20934 23738
rect 20804 23728 20934 23735
rect 21064 23735 21112 23848
rect 21146 23735 21194 23848
rect 21064 23728 21194 23735
rect 21324 23911 21454 23918
rect 21324 23798 21370 23911
rect 21404 23798 21454 23911
rect 21324 23738 21334 23798
rect 21444 23738 21454 23798
rect 21324 23735 21370 23738
rect 21404 23735 21454 23738
rect 21324 23728 21454 23735
rect 21574 23911 21704 23918
rect 21574 23908 21628 23911
rect 21662 23908 21704 23911
rect 21574 23848 21584 23908
rect 21694 23848 21704 23908
rect 21574 23735 21628 23848
rect 21662 23735 21704 23848
rect 21574 23728 21704 23735
rect 21844 23911 21974 23918
rect 21844 23798 21886 23911
rect 21920 23798 21974 23911
rect 21844 23738 21854 23798
rect 21964 23738 21974 23798
rect 21844 23735 21886 23738
rect 21920 23735 21974 23738
rect 21844 23728 21974 23735
rect 22094 23911 22224 23918
rect 22094 23908 22144 23911
rect 22178 23908 22224 23911
rect 22094 23848 22104 23908
rect 22214 23848 22224 23908
rect 22094 23735 22144 23848
rect 22178 23735 22224 23848
rect 22094 23728 22224 23735
rect 22354 23911 22484 23918
rect 22354 23798 22402 23911
rect 22436 23798 22484 23911
rect 22354 23738 22364 23798
rect 22474 23738 22484 23798
rect 22354 23735 22402 23738
rect 22436 23735 22484 23738
rect 22354 23728 22484 23735
rect 22614 23911 22744 23918
rect 22614 23908 22660 23911
rect 22694 23908 22744 23911
rect 22614 23848 22624 23908
rect 22734 23848 22744 23908
rect 22614 23735 22660 23848
rect 22694 23735 22744 23848
rect 22912 23911 22958 23923
rect 22912 23808 22918 23911
rect 22614 23728 22744 23735
rect 22864 23798 22918 23808
rect 22952 23808 22958 23911
rect 22994 23868 23004 24018
rect 23084 23868 23094 24018
rect 23170 23918 23216 23923
rect 22994 23838 23094 23868
rect 22952 23798 22994 23808
rect 22864 23738 22874 23798
rect 22984 23738 22994 23798
rect 22864 23735 22918 23738
rect 22952 23735 22994 23738
rect 22864 23728 22994 23735
rect 20590 23723 20636 23728
rect 20848 23723 20894 23728
rect 21106 23723 21152 23728
rect 21364 23723 21410 23728
rect 21622 23723 21668 23728
rect 21880 23723 21926 23728
rect 22138 23723 22184 23728
rect 22396 23723 22442 23728
rect 22654 23723 22700 23728
rect 22912 23723 22958 23728
rect 20334 23718 20384 23723
rect 20334 23691 20404 23718
rect 23024 23691 23094 23838
rect 23124 23911 23254 23918
rect 23124 23908 23176 23911
rect 23210 23908 23254 23911
rect 23124 23848 23134 23908
rect 23244 23848 23254 23908
rect 23124 23735 23176 23848
rect 23210 23735 23254 23848
rect 23124 23728 23254 23735
rect 23424 23911 23474 23928
rect 23424 23735 23434 23911
rect 23468 23735 23474 23911
rect 23170 23723 23216 23728
rect 23424 23718 23474 23735
rect 23394 23691 23474 23718
rect 20334 23688 20580 23691
rect 20334 23685 20584 23688
rect 20904 23685 21096 23691
rect 21162 23685 21354 23691
rect 21936 23685 22128 23691
rect 22194 23685 22386 23691
rect 22968 23685 23160 23691
rect 23226 23688 23474 23691
rect 23214 23685 23474 23688
rect 20334 23651 20400 23685
rect 20568 23651 20584 23685
rect 20900 23651 20916 23685
rect 21084 23651 21174 23685
rect 21342 23651 21948 23685
rect 22116 23651 22206 23685
rect 22374 23651 22980 23685
rect 23148 23651 23164 23685
rect 23214 23651 23238 23685
rect 23406 23651 23474 23685
rect 20334 23588 20584 23651
rect 20904 23645 21096 23651
rect 21162 23645 21354 23651
rect 21936 23645 22128 23651
rect 22194 23645 22386 23651
rect 22968 23645 23160 23651
rect 20334 23559 21104 23588
rect 21784 23578 21794 23608
rect 20334 23525 20400 23559
rect 20568 23525 20658 23559
rect 20826 23525 20916 23559
rect 21084 23525 21104 23559
rect 20334 23508 21104 23525
rect 21154 23559 21794 23578
rect 22014 23578 22024 23608
rect 23214 23588 23474 23651
rect 22014 23559 22654 23578
rect 21154 23525 21174 23559
rect 21342 23525 21432 23559
rect 21600 23525 21690 23559
rect 21858 23525 21948 23548
rect 22116 23525 22206 23559
rect 22374 23525 22464 23559
rect 22632 23525 22654 23559
rect 21154 23518 22654 23525
rect 22704 23559 23474 23588
rect 22704 23525 22722 23559
rect 22890 23525 22980 23559
rect 23148 23525 23238 23559
rect 23406 23525 23474 23559
rect 21784 23508 22024 23518
rect 20334 23488 21124 23508
rect 20334 23487 21148 23488
rect 20332 23475 21152 23487
rect 20332 23415 20338 23475
rect 20372 23415 20596 23475
rect 20630 23415 20854 23475
rect 20888 23415 21112 23475
rect 21146 23415 21152 23475
rect 20332 23403 21152 23415
rect 21344 23413 21359 23488
rect 21414 23413 21434 23488
rect 21344 23403 21434 23413
rect 21574 23475 21714 23488
rect 21574 23415 21628 23475
rect 21662 23415 21714 23475
rect 19738 23368 20224 23378
rect 19738 23248 19794 23368
rect 20214 23248 20224 23368
rect 19738 23238 20224 23248
rect 20334 23318 21148 23403
rect 21574 23318 21714 23415
rect 21859 23475 21949 23508
rect 22704 23488 23474 23525
rect 21859 23415 21886 23475
rect 21920 23415 21949 23475
rect 21859 23398 21949 23415
rect 22094 23475 22234 23488
rect 22094 23415 22144 23475
rect 22178 23415 22234 23475
rect 22094 23318 22234 23415
rect 22379 23413 22389 23488
rect 22444 23413 22454 23488
rect 22379 23403 22454 23413
rect 22654 23475 23474 23488
rect 22654 23415 22660 23475
rect 22694 23415 22918 23475
rect 22952 23415 23176 23475
rect 23210 23415 23434 23475
rect 23468 23415 23474 23475
rect 22654 23318 23474 23415
rect 20334 23298 23474 23318
rect 20334 23228 20354 23298
rect 23454 23228 23474 23298
rect 20334 23208 23474 23228
rect 23664 22938 23774 24738
rect 18864 22918 23774 22938
rect 18864 22868 20294 22918
rect 23504 22868 23774 22918
rect 23814 22828 23864 24848
rect 18764 22758 20294 22828
rect 23504 22758 23864 22828
rect 18764 22738 23864 22758
rect 23964 22638 24044 25038
rect 18604 22538 24044 22638
rect 24084 22498 24164 25178
rect 25684 25178 26304 25258
rect 25684 25078 25784 25178
rect 26204 25078 26304 25178
rect 26684 25078 27524 25118
rect 25544 25058 25804 25078
rect 24424 24898 24684 24918
rect 24424 24418 24444 24898
rect 24664 24418 24684 24898
rect 25544 24878 25564 25058
rect 25784 24878 25804 25058
rect 26184 25058 26444 25078
rect 25544 24867 25721 24878
rect 25755 24867 25804 24878
rect 25544 24858 25804 24867
rect 25973 25043 26019 25055
rect 25973 24867 25979 25043
rect 26013 24867 26019 25043
rect 25715 24855 25761 24858
rect 25973 24855 26019 24867
rect 26184 24878 26204 25058
rect 26424 24878 26444 25058
rect 26184 24867 26237 24878
rect 26271 24867 26444 24878
rect 26184 24858 26444 24867
rect 26484 25058 27224 25078
rect 26484 24878 26504 25058
rect 26604 24878 27224 25058
rect 26484 24858 27224 24878
rect 27304 24858 27524 25078
rect 26231 24855 26277 24858
rect 25771 24818 25963 24823
rect 26029 24818 26221 24823
rect 26684 24818 27524 24858
rect 25764 24817 26224 24818
rect 25764 24783 25783 24817
rect 25951 24783 26041 24817
rect 26209 24783 26224 24817
rect 25764 24718 26224 24783
rect 25764 24538 25784 24718
rect 26204 24538 26224 24718
rect 25764 24518 26224 24538
rect 24424 24398 24684 24418
rect 25764 24418 26224 24438
rect 25764 24238 25784 24418
rect 26204 24238 26224 24418
rect 25764 24172 26224 24238
rect 25764 24138 25783 24172
rect 25951 24138 26041 24172
rect 26209 24138 26224 24172
rect 25771 24132 25963 24138
rect 26029 24132 26221 24138
rect 26684 24098 27524 24138
rect 25544 24079 25804 24098
rect 25544 24078 25721 24079
rect 25755 24078 25804 24079
rect 25544 23898 25564 24078
rect 25784 23898 25804 24078
rect 25544 23878 25804 23898
rect 25944 24079 26044 24098
rect 25944 23903 25979 24079
rect 26013 23903 26044 24079
rect 25944 23798 26044 23903
rect 26184 24079 26444 24098
rect 26184 24078 26237 24079
rect 26271 24078 26444 24079
rect 26184 23898 26204 24078
rect 26424 23898 26444 24078
rect 26184 23878 26444 23898
rect 26484 24078 27524 24098
rect 26484 23898 26504 24078
rect 26604 23898 27404 24078
rect 26484 23878 27404 23898
rect 26684 23858 27404 23878
rect 27484 23858 27524 24078
rect 26684 23838 27524 23858
rect 25684 23718 26304 23798
rect 25684 23618 25784 23718
rect 26204 23618 26304 23718
rect 26684 23618 27524 23658
rect 25544 23598 25804 23618
rect 25544 23418 25564 23598
rect 25784 23418 25804 23598
rect 26184 23598 26444 23618
rect 25544 23407 25721 23418
rect 25755 23407 25804 23418
rect 25544 23398 25804 23407
rect 25973 23583 26019 23595
rect 25973 23407 25979 23583
rect 26013 23407 26019 23583
rect 25715 23395 25761 23398
rect 25973 23395 26019 23407
rect 26184 23418 26204 23598
rect 26424 23418 26444 23598
rect 26184 23407 26237 23418
rect 26271 23407 26444 23418
rect 26184 23398 26444 23407
rect 26484 23598 27224 23618
rect 26484 23418 26504 23598
rect 26604 23418 27224 23598
rect 26484 23398 27224 23418
rect 27304 23398 27524 23618
rect 26231 23395 26277 23398
rect 25771 23358 25963 23363
rect 26029 23358 26221 23363
rect 26684 23358 27524 23398
rect 25764 23357 26224 23358
rect 25764 23323 25783 23357
rect 25951 23323 26041 23357
rect 26209 23323 26224 23357
rect 24264 23298 24404 23318
rect 24264 22858 24284 23298
rect 24384 22858 24404 23298
rect 25764 23258 26224 23323
rect 25764 23078 25784 23258
rect 26204 23078 26224 23258
rect 25764 23058 26224 23078
rect 24264 22838 24404 22858
rect 25402 22718 26414 22738
rect 25402 22658 25424 22718
rect 26384 22707 26414 22718
rect 26385 22673 26414 22707
rect 26384 22658 26414 22673
rect 25402 22642 26414 22658
rect 18464 22438 24164 22498
rect 25044 22478 26044 22498
rect 24444 22439 24644 22458
rect 24444 22438 24486 22439
rect 24592 22438 24644 22439
rect 13436 22408 13836 22428
rect 12694 22308 13706 22324
rect 22364 22316 23524 22318
rect 12694 22248 12716 22308
rect 13696 22248 13706 22308
rect 12694 22228 13706 22248
rect 22360 22298 23524 22316
rect 10956 22088 11936 22108
rect 22360 22218 22384 22298
rect 23504 22218 23524 22298
rect 22360 22198 23524 22218
rect 22360 22146 22948 22198
rect 24444 22178 24464 22438
rect 22360 22040 22488 22146
rect 22885 22040 22948 22146
rect 22360 22004 22948 22040
rect 23664 22158 24464 22178
rect 23664 21978 23684 22158
rect 24624 21978 24644 22438
rect 25044 22298 25064 22478
rect 25244 22402 26044 22478
rect 25244 22368 25546 22402
rect 26034 22368 26044 22402
rect 25244 22298 26044 22368
rect 25044 22278 26044 22298
rect 26144 22478 26544 22498
rect 26144 22466 26344 22478
rect 26144 22302 26158 22466
rect 26206 22302 26344 22466
rect 26144 22298 26344 22302
rect 26524 22298 26544 22478
rect 26144 22278 26544 22298
rect 25402 22178 26414 22194
rect 25402 22118 25424 22178
rect 26404 22118 26414 22178
rect 25402 22098 26414 22118
rect 23664 21958 24644 21978
rect 12932 18962 13392 18982
rect 12932 18782 12952 18962
rect 13372 18782 13392 18962
rect 12932 18716 13392 18782
rect 12932 18682 12951 18716
rect 13119 18682 13209 18716
rect 13377 18682 13392 18716
rect 26114 18832 26574 18852
rect 12939 18676 13131 18682
rect 13197 18676 13389 18682
rect 13852 18642 14692 18682
rect 12712 18623 12972 18642
rect 12712 18622 12889 18623
rect 12923 18622 12972 18623
rect 12712 18442 12732 18622
rect 12952 18442 12972 18622
rect 12712 18422 12972 18442
rect 13112 18623 13212 18642
rect 13112 18447 13147 18623
rect 13181 18447 13212 18623
rect 13112 18342 13212 18447
rect 13352 18623 13612 18642
rect 13352 18622 13405 18623
rect 13439 18622 13612 18623
rect 13352 18442 13372 18622
rect 13592 18442 13612 18622
rect 13352 18422 13612 18442
rect 13652 18622 14692 18642
rect 13652 18442 13672 18622
rect 13772 18442 14572 18622
rect 13652 18422 14572 18442
rect 13852 18402 14572 18422
rect 14652 18402 14692 18622
rect 26114 18652 26134 18832
rect 26554 18652 26574 18832
rect 26114 18586 26574 18652
rect 26114 18552 26133 18586
rect 26301 18552 26391 18586
rect 26559 18552 26574 18586
rect 26121 18546 26313 18552
rect 26379 18546 26571 18552
rect 27034 18512 27874 18552
rect 13852 18382 14692 18402
rect 25894 18493 26154 18512
rect 25894 18492 26071 18493
rect 26105 18492 26154 18493
rect 5632 18302 11332 18322
rect 5632 18262 7462 18302
rect 10672 18262 11332 18302
rect 5632 15582 5732 18262
rect 5772 18142 7462 18222
rect 10672 18142 11212 18222
rect 5772 18122 11212 18142
rect 5772 15722 5832 18122
rect 5932 17932 11032 18022
rect 5932 15912 5992 17932
rect 6032 17822 10942 17892
rect 6032 16022 6132 17822
rect 6906 17582 10642 17602
rect 6906 17562 7462 17582
rect 6906 17522 7012 17562
rect 6906 17502 7462 17522
rect 10622 17502 10642 17582
rect 6906 17482 10642 17502
rect 7502 17434 7562 17482
rect 7500 17422 7562 17434
rect 7752 17432 7812 17442
rect 7500 17246 7506 17422
rect 7540 17246 7562 17422
rect 7500 17234 7562 17246
rect 7712 17422 7862 17432
rect 7712 17312 7764 17422
rect 7798 17312 7862 17422
rect 7712 17252 7722 17312
rect 7832 17252 7862 17312
rect 7712 17246 7764 17252
rect 7798 17246 7862 17252
rect 7712 17242 7862 17246
rect 7972 17422 8102 17482
rect 8274 17432 8320 17434
rect 7972 17246 8022 17422
rect 8056 17246 8102 17422
rect 7972 17242 8102 17246
rect 8232 17422 8362 17432
rect 8232 17312 8280 17422
rect 8314 17312 8362 17422
rect 8232 17252 8242 17312
rect 8352 17252 8362 17312
rect 8232 17246 8280 17252
rect 8314 17246 8362 17252
rect 8232 17242 8362 17246
rect 8492 17422 8622 17482
rect 8492 17246 8538 17422
rect 8572 17246 8622 17422
rect 8492 17242 8622 17246
rect 8742 17422 8872 17442
rect 8742 17312 8796 17422
rect 8830 17312 8872 17422
rect 7502 17193 7562 17234
rect 7752 17232 7862 17242
rect 8016 17234 8062 17242
rect 8274 17234 8320 17242
rect 8532 17234 8578 17242
rect 7812 17193 7862 17232
rect 8742 17202 8752 17312
rect 8862 17202 8872 17312
rect 9002 17422 9132 17482
rect 9306 17432 9352 17434
rect 9002 17246 9054 17422
rect 9088 17246 9132 17422
rect 9002 17242 9132 17246
rect 9262 17422 9392 17432
rect 9262 17322 9312 17422
rect 9346 17322 9392 17422
rect 9262 17252 9272 17322
rect 9382 17252 9392 17322
rect 9262 17246 9312 17252
rect 9346 17246 9392 17252
rect 9262 17242 9392 17246
rect 9522 17422 9652 17482
rect 9522 17246 9570 17422
rect 9604 17246 9652 17422
rect 9522 17242 9652 17246
rect 9782 17422 9912 17442
rect 9782 17322 9828 17422
rect 9862 17322 9912 17422
rect 9048 17234 9094 17242
rect 9306 17234 9352 17242
rect 9564 17234 9610 17242
rect 8742 17193 8872 17202
rect 9782 17202 9792 17322
rect 9902 17202 9912 17322
rect 10042 17422 10172 17482
rect 10602 17434 10642 17482
rect 10338 17432 10384 17434
rect 10042 17246 10086 17422
rect 10120 17246 10172 17422
rect 10042 17242 10172 17246
rect 10292 17422 10422 17432
rect 10292 17322 10344 17422
rect 10378 17322 10422 17422
rect 10292 17252 10302 17322
rect 10412 17252 10422 17322
rect 10292 17246 10344 17252
rect 10378 17246 10422 17252
rect 10292 17242 10422 17246
rect 10596 17422 10642 17434
rect 10596 17246 10602 17422
rect 10636 17246 10642 17422
rect 10080 17234 10126 17242
rect 10338 17234 10384 17242
rect 10596 17234 10642 17246
rect 10602 17202 10642 17234
rect 9782 17193 9912 17202
rect 7502 17192 7748 17193
rect 7502 17187 7752 17192
rect 7812 17187 8006 17193
rect 8072 17187 8264 17193
rect 8330 17187 8522 17193
rect 8588 17187 9038 17193
rect 9104 17187 9296 17193
rect 9362 17187 9554 17193
rect 9620 17187 10070 17193
rect 10136 17187 10328 17193
rect 10392 17187 10642 17202
rect 7502 17153 7568 17187
rect 7736 17153 7752 17187
rect 7810 17153 7826 17187
rect 7994 17153 8084 17187
rect 8252 17153 8342 17187
rect 8510 17153 8600 17187
rect 8768 17153 8858 17187
rect 9026 17153 9116 17187
rect 9284 17153 9374 17187
rect 9542 17153 9632 17187
rect 9800 17153 9890 17187
rect 10058 17153 10148 17187
rect 10316 17153 10332 17187
rect 10392 17153 10406 17187
rect 10574 17153 10642 17187
rect 7502 17152 7752 17153
rect 7812 17152 8006 17153
rect 7556 17147 7748 17152
rect 7814 17147 8006 17152
rect 8072 17147 8264 17153
rect 8330 17147 8522 17153
rect 8588 17147 8780 17153
rect 8846 17147 9038 17153
rect 9104 17147 9296 17153
rect 9362 17147 9554 17153
rect 9620 17147 9812 17153
rect 9878 17147 10070 17153
rect 10136 17147 10328 17153
rect 10392 17152 10642 17153
rect 10394 17147 10586 17152
rect 8092 17102 8202 17112
rect 7814 17079 8006 17085
rect 8092 17079 8102 17102
rect 7810 17045 7826 17079
rect 7994 17045 8102 17079
rect 7814 17039 8006 17045
rect 7502 17007 7552 17012
rect 7500 16995 7552 17007
rect 7758 17002 7804 17007
rect 7500 16819 7506 16995
rect 7540 16819 7552 16995
rect 7500 16807 7552 16819
rect 7712 16995 7842 17002
rect 7712 16992 7764 16995
rect 7798 16992 7842 16995
rect 7712 16932 7722 16992
rect 7832 16932 7842 16992
rect 7712 16819 7764 16932
rect 7798 16819 7842 16932
rect 8016 16995 8062 17007
rect 8016 16902 8022 16995
rect 7712 16812 7842 16819
rect 7972 16882 8022 16902
rect 8056 16902 8062 16995
rect 8092 16942 8102 17045
rect 8192 17079 8202 17102
rect 10162 17102 10262 17112
rect 8588 17079 8780 17085
rect 8846 17079 9038 17085
rect 9620 17079 9812 17085
rect 9878 17079 10070 17085
rect 8192 17045 8600 17079
rect 8768 17045 8858 17079
rect 9026 17045 9632 17079
rect 9800 17045 9890 17079
rect 10058 17045 10074 17079
rect 8192 16942 8202 17045
rect 8588 17039 8780 17045
rect 8846 17039 9038 17045
rect 9620 17039 9812 17045
rect 9878 17039 10070 17045
rect 8274 17002 8320 17007
rect 8532 17002 8578 17007
rect 8790 17002 8836 17007
rect 9048 17002 9094 17007
rect 9306 17002 9352 17007
rect 9564 17002 9610 17007
rect 9822 17002 9868 17007
rect 8092 16932 8202 16942
rect 8232 16995 8362 17002
rect 8232 16992 8280 16995
rect 8314 16992 8362 16995
rect 8232 16932 8242 16992
rect 8352 16932 8362 16992
rect 8056 16882 8102 16902
rect 7972 16822 7982 16882
rect 8092 16822 8102 16882
rect 7972 16819 8022 16822
rect 8056 16819 8102 16822
rect 7972 16812 8102 16819
rect 8232 16819 8280 16932
rect 8314 16819 8362 16932
rect 8232 16812 8362 16819
rect 8492 16995 8622 17002
rect 8492 16882 8538 16995
rect 8572 16882 8622 16995
rect 8492 16822 8502 16882
rect 8612 16822 8622 16882
rect 8492 16819 8538 16822
rect 8572 16819 8622 16822
rect 8492 16812 8622 16819
rect 8742 16995 8872 17002
rect 8742 16992 8796 16995
rect 8830 16992 8872 16995
rect 8742 16932 8752 16992
rect 8862 16932 8872 16992
rect 8742 16819 8796 16932
rect 8830 16819 8872 16932
rect 8742 16812 8872 16819
rect 9012 16995 9142 17002
rect 9012 16882 9054 16995
rect 9088 16882 9142 16995
rect 9012 16822 9022 16882
rect 9132 16822 9142 16882
rect 9012 16819 9054 16822
rect 9088 16819 9142 16822
rect 9012 16812 9142 16819
rect 9262 16995 9392 17002
rect 9262 16992 9312 16995
rect 9346 16992 9392 16995
rect 9262 16932 9272 16992
rect 9382 16932 9392 16992
rect 9262 16819 9312 16932
rect 9346 16819 9392 16932
rect 9262 16812 9392 16819
rect 9522 16995 9652 17002
rect 9522 16882 9570 16995
rect 9604 16882 9652 16995
rect 9522 16822 9532 16882
rect 9642 16822 9652 16882
rect 9522 16819 9570 16822
rect 9604 16819 9652 16822
rect 9522 16812 9652 16819
rect 9782 16995 9912 17002
rect 9782 16992 9828 16995
rect 9862 16992 9912 16995
rect 9782 16932 9792 16992
rect 9902 16932 9912 16992
rect 9782 16819 9828 16932
rect 9862 16819 9912 16932
rect 10080 16995 10126 17007
rect 10080 16892 10086 16995
rect 9782 16812 9912 16819
rect 10032 16882 10086 16892
rect 10120 16892 10126 16995
rect 10162 16952 10172 17102
rect 10252 16952 10262 17102
rect 10338 17002 10384 17007
rect 10162 16922 10262 16952
rect 10120 16882 10162 16892
rect 10032 16822 10042 16882
rect 10152 16822 10162 16882
rect 10032 16819 10086 16822
rect 10120 16819 10162 16822
rect 10032 16812 10162 16819
rect 7758 16807 7804 16812
rect 8016 16807 8062 16812
rect 8274 16807 8320 16812
rect 8532 16807 8578 16812
rect 8790 16807 8836 16812
rect 9048 16807 9094 16812
rect 9306 16807 9352 16812
rect 9564 16807 9610 16812
rect 9822 16807 9868 16812
rect 10080 16807 10126 16812
rect 7502 16802 7552 16807
rect 7502 16775 7572 16802
rect 10192 16775 10262 16922
rect 10292 16995 10422 17002
rect 10292 16992 10344 16995
rect 10378 16992 10422 16995
rect 10292 16932 10302 16992
rect 10412 16932 10422 16992
rect 10292 16819 10344 16932
rect 10378 16819 10422 16932
rect 10292 16812 10422 16819
rect 10592 16995 10642 17012
rect 10592 16819 10602 16995
rect 10636 16819 10642 16995
rect 10338 16807 10384 16812
rect 10592 16802 10642 16819
rect 10562 16775 10642 16802
rect 7502 16772 7748 16775
rect 7502 16769 7752 16772
rect 8072 16769 8264 16775
rect 8330 16769 8522 16775
rect 9104 16769 9296 16775
rect 9362 16769 9554 16775
rect 10136 16769 10328 16775
rect 10394 16772 10642 16775
rect 10382 16769 10642 16772
rect 7502 16735 7568 16769
rect 7736 16735 7752 16769
rect 8068 16735 8084 16769
rect 8252 16735 8342 16769
rect 8510 16735 9116 16769
rect 9284 16735 9374 16769
rect 9542 16735 10148 16769
rect 10316 16735 10332 16769
rect 10382 16735 10406 16769
rect 10574 16735 10642 16769
rect 7502 16672 7752 16735
rect 8072 16729 8264 16735
rect 8330 16729 8522 16735
rect 9104 16729 9296 16735
rect 9362 16729 9554 16735
rect 10136 16729 10328 16735
rect 7502 16643 8272 16672
rect 8952 16662 8962 16692
rect 7502 16609 7568 16643
rect 7736 16609 7826 16643
rect 7994 16609 8084 16643
rect 8252 16609 8272 16643
rect 7502 16592 8272 16609
rect 8322 16643 8962 16662
rect 9182 16662 9192 16692
rect 10382 16672 10642 16735
rect 9182 16643 9822 16662
rect 8322 16609 8342 16643
rect 8510 16609 8600 16643
rect 8768 16609 8858 16643
rect 9026 16609 9116 16632
rect 9284 16609 9374 16643
rect 9542 16609 9632 16643
rect 9800 16609 9822 16643
rect 8322 16602 9822 16609
rect 9872 16643 10642 16672
rect 9872 16609 9890 16643
rect 10058 16609 10148 16643
rect 10316 16609 10406 16643
rect 10574 16609 10642 16643
rect 8952 16592 9192 16602
rect 7502 16572 8292 16592
rect 7502 16571 8316 16572
rect 7500 16559 8320 16571
rect 7500 16499 7506 16559
rect 7540 16499 7764 16559
rect 7798 16499 8022 16559
rect 8056 16499 8280 16559
rect 8314 16499 8320 16559
rect 7500 16487 8320 16499
rect 8512 16497 8527 16572
rect 8582 16497 8602 16572
rect 8512 16487 8602 16497
rect 8742 16559 8882 16572
rect 8742 16499 8796 16559
rect 8830 16499 8882 16559
rect 6906 16452 7392 16462
rect 6906 16332 6962 16452
rect 7382 16332 7392 16452
rect 6906 16322 7392 16332
rect 7502 16402 8316 16487
rect 8742 16402 8882 16499
rect 9027 16559 9117 16592
rect 9872 16572 10642 16609
rect 9027 16499 9054 16559
rect 9088 16499 9117 16559
rect 9027 16482 9117 16499
rect 9262 16559 9402 16572
rect 9262 16499 9312 16559
rect 9346 16499 9402 16559
rect 9262 16402 9402 16499
rect 9547 16497 9557 16572
rect 9612 16497 9622 16572
rect 9547 16487 9622 16497
rect 9822 16559 10642 16572
rect 9822 16499 9828 16559
rect 9862 16499 10086 16559
rect 10120 16499 10344 16559
rect 10378 16499 10602 16559
rect 10636 16499 10642 16559
rect 9822 16402 10642 16499
rect 7502 16382 10642 16402
rect 7502 16312 7522 16382
rect 10622 16312 10642 16382
rect 7502 16292 10642 16312
rect 10832 16022 10942 17822
rect 6032 16002 10942 16022
rect 6032 15952 7462 16002
rect 10672 15952 10942 16002
rect 10982 15912 11032 17932
rect 5932 15842 7462 15912
rect 10672 15842 11032 15912
rect 5932 15822 11032 15842
rect 11132 15722 11212 18122
rect 5772 15622 11212 15722
rect 11252 15582 11332 18262
rect 12852 18262 13472 18342
rect 25894 18312 25914 18492
rect 26134 18312 26154 18492
rect 25894 18292 26154 18312
rect 26294 18493 26394 18512
rect 26294 18317 26329 18493
rect 26363 18317 26394 18493
rect 12852 18162 12952 18262
rect 13372 18162 13472 18262
rect 26294 18212 26394 18317
rect 26534 18493 26794 18512
rect 26534 18492 26587 18493
rect 26621 18492 26794 18493
rect 26534 18312 26554 18492
rect 26774 18312 26794 18492
rect 26534 18292 26794 18312
rect 26834 18492 27874 18512
rect 26834 18312 26854 18492
rect 26954 18312 27754 18492
rect 26834 18292 27754 18312
rect 27034 18272 27754 18292
rect 27834 18272 27874 18492
rect 27034 18252 27874 18272
rect 13852 18162 14692 18202
rect 12712 18142 12972 18162
rect 11592 17982 11852 18002
rect 11592 17502 11612 17982
rect 11832 17502 11852 17982
rect 12712 17962 12732 18142
rect 12952 17962 12972 18142
rect 13352 18142 13612 18162
rect 12712 17951 12889 17962
rect 12923 17951 12972 17962
rect 12712 17942 12972 17951
rect 13141 18127 13187 18139
rect 13141 17951 13147 18127
rect 13181 17951 13187 18127
rect 12883 17939 12929 17942
rect 13141 17939 13187 17951
rect 13352 17962 13372 18142
rect 13592 17962 13612 18142
rect 13352 17951 13405 17962
rect 13439 17951 13612 17962
rect 13352 17942 13612 17951
rect 13652 18142 14392 18162
rect 13652 17962 13672 18142
rect 13772 17962 14392 18142
rect 13652 17942 14392 17962
rect 14472 17942 14692 18162
rect 13399 17939 13445 17942
rect 12939 17902 13131 17907
rect 13197 17902 13389 17907
rect 13852 17902 14692 17942
rect 18814 18172 24514 18192
rect 18814 18132 20644 18172
rect 23854 18132 24514 18172
rect 12932 17901 13392 17902
rect 12932 17867 12951 17901
rect 13119 17867 13209 17901
rect 13377 17867 13392 17901
rect 12932 17802 13392 17867
rect 12932 17622 12952 17802
rect 13372 17622 13392 17802
rect 12932 17602 13392 17622
rect 11592 17482 11852 17502
rect 12932 17502 13392 17522
rect 12932 17322 12952 17502
rect 13372 17322 13392 17502
rect 12932 17256 13392 17322
rect 12932 17222 12951 17256
rect 13119 17222 13209 17256
rect 13377 17222 13392 17256
rect 12939 17216 13131 17222
rect 13197 17216 13389 17222
rect 13852 17182 14692 17222
rect 12712 17163 12972 17182
rect 12712 17162 12889 17163
rect 12923 17162 12972 17163
rect 12712 16982 12732 17162
rect 12952 16982 12972 17162
rect 12712 16962 12972 16982
rect 13112 17163 13212 17182
rect 13112 16987 13147 17163
rect 13181 16987 13212 17163
rect 13112 16882 13212 16987
rect 13352 17163 13612 17182
rect 13352 17162 13405 17163
rect 13439 17162 13612 17163
rect 13352 16982 13372 17162
rect 13592 16982 13612 17162
rect 13352 16962 13612 16982
rect 13652 17162 14692 17182
rect 13652 16982 13672 17162
rect 13772 16982 14572 17162
rect 13652 16962 14572 16982
rect 13852 16942 14572 16962
rect 14652 16942 14692 17162
rect 13852 16922 14692 16942
rect 12852 16802 13472 16882
rect 12852 16702 12952 16802
rect 13372 16702 13472 16802
rect 13852 16702 14692 16742
rect 12712 16682 12972 16702
rect 12712 16502 12732 16682
rect 12952 16502 12972 16682
rect 13352 16682 13612 16702
rect 12712 16491 12889 16502
rect 12923 16491 12972 16502
rect 12712 16482 12972 16491
rect 13141 16667 13187 16679
rect 13141 16491 13147 16667
rect 13181 16491 13187 16667
rect 12883 16479 12929 16482
rect 13141 16479 13187 16491
rect 13352 16502 13372 16682
rect 13592 16502 13612 16682
rect 13352 16491 13405 16502
rect 13439 16491 13612 16502
rect 13352 16482 13612 16491
rect 13652 16682 14392 16702
rect 13652 16502 13672 16682
rect 13772 16502 14392 16682
rect 13652 16482 14392 16502
rect 14472 16482 14692 16702
rect 13399 16479 13445 16482
rect 12939 16442 13131 16447
rect 13197 16442 13389 16447
rect 13852 16442 14692 16482
rect 12932 16441 13392 16442
rect 12932 16407 12951 16441
rect 13119 16407 13209 16441
rect 13377 16407 13392 16441
rect 11432 16382 11572 16402
rect 11432 15942 11452 16382
rect 11552 15942 11572 16382
rect 12932 16342 13392 16407
rect 12932 16162 12952 16342
rect 13372 16162 13392 16342
rect 12932 16142 13392 16162
rect 11432 15922 11572 15942
rect 12570 15802 13582 15822
rect 12570 15742 12592 15802
rect 13552 15791 13582 15802
rect 13553 15757 13582 15791
rect 13552 15742 13582 15757
rect 12570 15726 13582 15742
rect 5632 15522 11332 15582
rect 12212 15562 13212 15582
rect 11612 15523 11812 15542
rect 11612 15522 11654 15523
rect 11760 15522 11812 15523
rect 9532 15400 10692 15402
rect 9528 15382 10692 15400
rect 9528 15302 9552 15382
rect 10672 15302 10692 15382
rect 9528 15282 10692 15302
rect 9528 15230 10116 15282
rect 11612 15262 11632 15522
rect 9528 15124 9656 15230
rect 10053 15124 10116 15230
rect 9528 15088 10116 15124
rect 10832 15242 11632 15262
rect 10832 15062 10852 15242
rect 11792 15062 11812 15522
rect 12212 15382 12232 15562
rect 12412 15486 13212 15562
rect 12412 15452 12714 15486
rect 13202 15452 13212 15486
rect 12412 15382 13212 15452
rect 12212 15362 13212 15382
rect 13312 15562 13712 15582
rect 13312 15550 13512 15562
rect 13312 15386 13326 15550
rect 13374 15386 13512 15550
rect 13312 15382 13512 15386
rect 13692 15382 13712 15562
rect 18814 15452 18914 18132
rect 18954 18012 20644 18092
rect 23854 18012 24394 18092
rect 18954 17992 24394 18012
rect 18954 15592 19014 17992
rect 19114 17802 24214 17892
rect 19114 15782 19174 17802
rect 19214 17692 24124 17762
rect 19214 15892 19314 17692
rect 20088 17452 23824 17472
rect 20088 17432 20644 17452
rect 20088 17392 20194 17432
rect 20088 17372 20644 17392
rect 23804 17372 23824 17452
rect 20088 17352 23824 17372
rect 20684 17304 20744 17352
rect 20682 17292 20744 17304
rect 20934 17302 20994 17312
rect 20682 17116 20688 17292
rect 20722 17116 20744 17292
rect 20682 17104 20744 17116
rect 20894 17292 21044 17302
rect 20894 17182 20946 17292
rect 20980 17182 21044 17292
rect 20894 17122 20904 17182
rect 21014 17122 21044 17182
rect 20894 17116 20946 17122
rect 20980 17116 21044 17122
rect 20894 17112 21044 17116
rect 21154 17292 21284 17352
rect 21456 17302 21502 17304
rect 21154 17116 21204 17292
rect 21238 17116 21284 17292
rect 21154 17112 21284 17116
rect 21414 17292 21544 17302
rect 21414 17182 21462 17292
rect 21496 17182 21544 17292
rect 21414 17122 21424 17182
rect 21534 17122 21544 17182
rect 21414 17116 21462 17122
rect 21496 17116 21544 17122
rect 21414 17112 21544 17116
rect 21674 17292 21804 17352
rect 21674 17116 21720 17292
rect 21754 17116 21804 17292
rect 21674 17112 21804 17116
rect 21924 17292 22054 17312
rect 21924 17182 21978 17292
rect 22012 17182 22054 17292
rect 20684 17063 20744 17104
rect 20934 17102 21044 17112
rect 21198 17104 21244 17112
rect 21456 17104 21502 17112
rect 21714 17104 21760 17112
rect 20994 17063 21044 17102
rect 21924 17072 21934 17182
rect 22044 17072 22054 17182
rect 22184 17292 22314 17352
rect 22488 17302 22534 17304
rect 22184 17116 22236 17292
rect 22270 17116 22314 17292
rect 22184 17112 22314 17116
rect 22444 17292 22574 17302
rect 22444 17192 22494 17292
rect 22528 17192 22574 17292
rect 22444 17122 22454 17192
rect 22564 17122 22574 17192
rect 22444 17116 22494 17122
rect 22528 17116 22574 17122
rect 22444 17112 22574 17116
rect 22704 17292 22834 17352
rect 22704 17116 22752 17292
rect 22786 17116 22834 17292
rect 22704 17112 22834 17116
rect 22964 17292 23094 17312
rect 22964 17192 23010 17292
rect 23044 17192 23094 17292
rect 22230 17104 22276 17112
rect 22488 17104 22534 17112
rect 22746 17104 22792 17112
rect 21924 17063 22054 17072
rect 22964 17072 22974 17192
rect 23084 17072 23094 17192
rect 23224 17292 23354 17352
rect 23784 17304 23824 17352
rect 23520 17302 23566 17304
rect 23224 17116 23268 17292
rect 23302 17116 23354 17292
rect 23224 17112 23354 17116
rect 23474 17292 23604 17302
rect 23474 17192 23526 17292
rect 23560 17192 23604 17292
rect 23474 17122 23484 17192
rect 23594 17122 23604 17192
rect 23474 17116 23526 17122
rect 23560 17116 23604 17122
rect 23474 17112 23604 17116
rect 23778 17292 23824 17304
rect 23778 17116 23784 17292
rect 23818 17116 23824 17292
rect 23262 17104 23308 17112
rect 23520 17104 23566 17112
rect 23778 17104 23824 17116
rect 23784 17072 23824 17104
rect 22964 17063 23094 17072
rect 20684 17062 20930 17063
rect 20684 17057 20934 17062
rect 20994 17057 21188 17063
rect 21254 17057 21446 17063
rect 21512 17057 21704 17063
rect 21770 17057 22220 17063
rect 22286 17057 22478 17063
rect 22544 17057 22736 17063
rect 22802 17057 23252 17063
rect 23318 17057 23510 17063
rect 23574 17057 23824 17072
rect 20684 17023 20750 17057
rect 20918 17023 20934 17057
rect 20992 17023 21008 17057
rect 21176 17023 21266 17057
rect 21434 17023 21524 17057
rect 21692 17023 21782 17057
rect 21950 17023 22040 17057
rect 22208 17023 22298 17057
rect 22466 17023 22556 17057
rect 22724 17023 22814 17057
rect 22982 17023 23072 17057
rect 23240 17023 23330 17057
rect 23498 17023 23514 17057
rect 23574 17023 23588 17057
rect 23756 17023 23824 17057
rect 20684 17022 20934 17023
rect 20994 17022 21188 17023
rect 20738 17017 20930 17022
rect 20996 17017 21188 17022
rect 21254 17017 21446 17023
rect 21512 17017 21704 17023
rect 21770 17017 21962 17023
rect 22028 17017 22220 17023
rect 22286 17017 22478 17023
rect 22544 17017 22736 17023
rect 22802 17017 22994 17023
rect 23060 17017 23252 17023
rect 23318 17017 23510 17023
rect 23574 17022 23824 17023
rect 23576 17017 23768 17022
rect 21274 16972 21384 16982
rect 20996 16949 21188 16955
rect 21274 16949 21284 16972
rect 20992 16915 21008 16949
rect 21176 16915 21284 16949
rect 20996 16909 21188 16915
rect 20684 16877 20734 16882
rect 20682 16865 20734 16877
rect 20940 16872 20986 16877
rect 20682 16689 20688 16865
rect 20722 16689 20734 16865
rect 20682 16677 20734 16689
rect 20894 16865 21024 16872
rect 20894 16862 20946 16865
rect 20980 16862 21024 16865
rect 20894 16802 20904 16862
rect 21014 16802 21024 16862
rect 20894 16689 20946 16802
rect 20980 16689 21024 16802
rect 21198 16865 21244 16877
rect 21198 16772 21204 16865
rect 20894 16682 21024 16689
rect 21154 16752 21204 16772
rect 21238 16772 21244 16865
rect 21274 16812 21284 16915
rect 21374 16949 21384 16972
rect 23344 16972 23444 16982
rect 21770 16949 21962 16955
rect 22028 16949 22220 16955
rect 22802 16949 22994 16955
rect 23060 16949 23252 16955
rect 21374 16915 21782 16949
rect 21950 16915 22040 16949
rect 22208 16915 22814 16949
rect 22982 16915 23072 16949
rect 23240 16915 23256 16949
rect 21374 16812 21384 16915
rect 21770 16909 21962 16915
rect 22028 16909 22220 16915
rect 22802 16909 22994 16915
rect 23060 16909 23252 16915
rect 21456 16872 21502 16877
rect 21714 16872 21760 16877
rect 21972 16872 22018 16877
rect 22230 16872 22276 16877
rect 22488 16872 22534 16877
rect 22746 16872 22792 16877
rect 23004 16872 23050 16877
rect 21274 16802 21384 16812
rect 21414 16865 21544 16872
rect 21414 16862 21462 16865
rect 21496 16862 21544 16865
rect 21414 16802 21424 16862
rect 21534 16802 21544 16862
rect 21238 16752 21284 16772
rect 21154 16692 21164 16752
rect 21274 16692 21284 16752
rect 21154 16689 21204 16692
rect 21238 16689 21284 16692
rect 21154 16682 21284 16689
rect 21414 16689 21462 16802
rect 21496 16689 21544 16802
rect 21414 16682 21544 16689
rect 21674 16865 21804 16872
rect 21674 16752 21720 16865
rect 21754 16752 21804 16865
rect 21674 16692 21684 16752
rect 21794 16692 21804 16752
rect 21674 16689 21720 16692
rect 21754 16689 21804 16692
rect 21674 16682 21804 16689
rect 21924 16865 22054 16872
rect 21924 16862 21978 16865
rect 22012 16862 22054 16865
rect 21924 16802 21934 16862
rect 22044 16802 22054 16862
rect 21924 16689 21978 16802
rect 22012 16689 22054 16802
rect 21924 16682 22054 16689
rect 22194 16865 22324 16872
rect 22194 16752 22236 16865
rect 22270 16752 22324 16865
rect 22194 16692 22204 16752
rect 22314 16692 22324 16752
rect 22194 16689 22236 16692
rect 22270 16689 22324 16692
rect 22194 16682 22324 16689
rect 22444 16865 22574 16872
rect 22444 16862 22494 16865
rect 22528 16862 22574 16865
rect 22444 16802 22454 16862
rect 22564 16802 22574 16862
rect 22444 16689 22494 16802
rect 22528 16689 22574 16802
rect 22444 16682 22574 16689
rect 22704 16865 22834 16872
rect 22704 16752 22752 16865
rect 22786 16752 22834 16865
rect 22704 16692 22714 16752
rect 22824 16692 22834 16752
rect 22704 16689 22752 16692
rect 22786 16689 22834 16692
rect 22704 16682 22834 16689
rect 22964 16865 23094 16872
rect 22964 16862 23010 16865
rect 23044 16862 23094 16865
rect 22964 16802 22974 16862
rect 23084 16802 23094 16862
rect 22964 16689 23010 16802
rect 23044 16689 23094 16802
rect 23262 16865 23308 16877
rect 23262 16762 23268 16865
rect 22964 16682 23094 16689
rect 23214 16752 23268 16762
rect 23302 16762 23308 16865
rect 23344 16822 23354 16972
rect 23434 16822 23444 16972
rect 23520 16872 23566 16877
rect 23344 16792 23444 16822
rect 23302 16752 23344 16762
rect 23214 16692 23224 16752
rect 23334 16692 23344 16752
rect 23214 16689 23268 16692
rect 23302 16689 23344 16692
rect 23214 16682 23344 16689
rect 20940 16677 20986 16682
rect 21198 16677 21244 16682
rect 21456 16677 21502 16682
rect 21714 16677 21760 16682
rect 21972 16677 22018 16682
rect 22230 16677 22276 16682
rect 22488 16677 22534 16682
rect 22746 16677 22792 16682
rect 23004 16677 23050 16682
rect 23262 16677 23308 16682
rect 20684 16672 20734 16677
rect 20684 16645 20754 16672
rect 23374 16645 23444 16792
rect 23474 16865 23604 16872
rect 23474 16862 23526 16865
rect 23560 16862 23604 16865
rect 23474 16802 23484 16862
rect 23594 16802 23604 16862
rect 23474 16689 23526 16802
rect 23560 16689 23604 16802
rect 23474 16682 23604 16689
rect 23774 16865 23824 16882
rect 23774 16689 23784 16865
rect 23818 16689 23824 16865
rect 23520 16677 23566 16682
rect 23774 16672 23824 16689
rect 23744 16645 23824 16672
rect 20684 16642 20930 16645
rect 20684 16639 20934 16642
rect 21254 16639 21446 16645
rect 21512 16639 21704 16645
rect 22286 16639 22478 16645
rect 22544 16639 22736 16645
rect 23318 16639 23510 16645
rect 23576 16642 23824 16645
rect 23564 16639 23824 16642
rect 20684 16605 20750 16639
rect 20918 16605 20934 16639
rect 21250 16605 21266 16639
rect 21434 16605 21524 16639
rect 21692 16605 22298 16639
rect 22466 16605 22556 16639
rect 22724 16605 23330 16639
rect 23498 16605 23514 16639
rect 23564 16605 23588 16639
rect 23756 16605 23824 16639
rect 20684 16542 20934 16605
rect 21254 16599 21446 16605
rect 21512 16599 21704 16605
rect 22286 16599 22478 16605
rect 22544 16599 22736 16605
rect 23318 16599 23510 16605
rect 20684 16513 21454 16542
rect 22134 16532 22144 16562
rect 20684 16479 20750 16513
rect 20918 16479 21008 16513
rect 21176 16479 21266 16513
rect 21434 16479 21454 16513
rect 20684 16462 21454 16479
rect 21504 16513 22144 16532
rect 22364 16532 22374 16562
rect 23564 16542 23824 16605
rect 22364 16513 23004 16532
rect 21504 16479 21524 16513
rect 21692 16479 21782 16513
rect 21950 16479 22040 16513
rect 22208 16479 22298 16502
rect 22466 16479 22556 16513
rect 22724 16479 22814 16513
rect 22982 16479 23004 16513
rect 21504 16472 23004 16479
rect 23054 16513 23824 16542
rect 23054 16479 23072 16513
rect 23240 16479 23330 16513
rect 23498 16479 23588 16513
rect 23756 16479 23824 16513
rect 22134 16462 22374 16472
rect 20684 16442 21474 16462
rect 20684 16441 21498 16442
rect 20682 16429 21502 16441
rect 20682 16369 20688 16429
rect 20722 16369 20946 16429
rect 20980 16369 21204 16429
rect 21238 16369 21462 16429
rect 21496 16369 21502 16429
rect 20682 16357 21502 16369
rect 21694 16367 21709 16442
rect 21764 16367 21784 16442
rect 21694 16357 21784 16367
rect 21924 16429 22064 16442
rect 21924 16369 21978 16429
rect 22012 16369 22064 16429
rect 20088 16322 20574 16332
rect 20088 16202 20144 16322
rect 20564 16202 20574 16322
rect 20088 16192 20574 16202
rect 20684 16272 21498 16357
rect 21924 16272 22064 16369
rect 22209 16429 22299 16462
rect 23054 16442 23824 16479
rect 22209 16369 22236 16429
rect 22270 16369 22299 16429
rect 22209 16352 22299 16369
rect 22444 16429 22584 16442
rect 22444 16369 22494 16429
rect 22528 16369 22584 16429
rect 22444 16272 22584 16369
rect 22729 16367 22739 16442
rect 22794 16367 22804 16442
rect 22729 16357 22804 16367
rect 23004 16429 23824 16442
rect 23004 16369 23010 16429
rect 23044 16369 23268 16429
rect 23302 16369 23526 16429
rect 23560 16369 23784 16429
rect 23818 16369 23824 16429
rect 23004 16272 23824 16369
rect 20684 16252 23824 16272
rect 20684 16182 20704 16252
rect 23804 16182 23824 16252
rect 20684 16162 23824 16182
rect 24014 15892 24124 17692
rect 19214 15872 24124 15892
rect 19214 15822 20644 15872
rect 23854 15822 24124 15872
rect 24164 15782 24214 17802
rect 19114 15712 20644 15782
rect 23854 15712 24214 15782
rect 19114 15692 24214 15712
rect 24314 15592 24394 17992
rect 18954 15492 24394 15592
rect 24434 15452 24514 18132
rect 26034 18132 26654 18212
rect 26034 18032 26134 18132
rect 26554 18032 26654 18132
rect 27034 18032 27874 18072
rect 25894 18012 26154 18032
rect 24774 17852 25034 17872
rect 24774 17372 24794 17852
rect 25014 17372 25034 17852
rect 25894 17832 25914 18012
rect 26134 17832 26154 18012
rect 26534 18012 26794 18032
rect 25894 17821 26071 17832
rect 26105 17821 26154 17832
rect 25894 17812 26154 17821
rect 26323 17997 26369 18009
rect 26323 17821 26329 17997
rect 26363 17821 26369 17997
rect 26065 17809 26111 17812
rect 26323 17809 26369 17821
rect 26534 17832 26554 18012
rect 26774 17832 26794 18012
rect 26534 17821 26587 17832
rect 26621 17821 26794 17832
rect 26534 17812 26794 17821
rect 26834 18012 27574 18032
rect 26834 17832 26854 18012
rect 26954 17832 27574 18012
rect 26834 17812 27574 17832
rect 27654 17812 27874 18032
rect 26581 17809 26627 17812
rect 26121 17772 26313 17777
rect 26379 17772 26571 17777
rect 27034 17772 27874 17812
rect 26114 17771 26574 17772
rect 26114 17737 26133 17771
rect 26301 17737 26391 17771
rect 26559 17737 26574 17771
rect 26114 17672 26574 17737
rect 26114 17492 26134 17672
rect 26554 17492 26574 17672
rect 26114 17472 26574 17492
rect 24774 17352 25034 17372
rect 26114 17372 26574 17392
rect 26114 17192 26134 17372
rect 26554 17192 26574 17372
rect 26114 17126 26574 17192
rect 26114 17092 26133 17126
rect 26301 17092 26391 17126
rect 26559 17092 26574 17126
rect 26121 17086 26313 17092
rect 26379 17086 26571 17092
rect 27034 17052 27874 17092
rect 25894 17033 26154 17052
rect 25894 17032 26071 17033
rect 26105 17032 26154 17033
rect 25894 16852 25914 17032
rect 26134 16852 26154 17032
rect 25894 16832 26154 16852
rect 26294 17033 26394 17052
rect 26294 16857 26329 17033
rect 26363 16857 26394 17033
rect 26294 16752 26394 16857
rect 26534 17033 26794 17052
rect 26534 17032 26587 17033
rect 26621 17032 26794 17033
rect 26534 16852 26554 17032
rect 26774 16852 26794 17032
rect 26534 16832 26794 16852
rect 26834 17032 27874 17052
rect 26834 16852 26854 17032
rect 26954 16852 27754 17032
rect 26834 16832 27754 16852
rect 27034 16812 27754 16832
rect 27834 16812 27874 17032
rect 27034 16792 27874 16812
rect 26034 16672 26654 16752
rect 26034 16572 26134 16672
rect 26554 16572 26654 16672
rect 27034 16572 27874 16612
rect 25894 16552 26154 16572
rect 25894 16372 25914 16552
rect 26134 16372 26154 16552
rect 26534 16552 26794 16572
rect 25894 16361 26071 16372
rect 26105 16361 26154 16372
rect 25894 16352 26154 16361
rect 26323 16537 26369 16549
rect 26323 16361 26329 16537
rect 26363 16361 26369 16537
rect 26065 16349 26111 16352
rect 26323 16349 26369 16361
rect 26534 16372 26554 16552
rect 26774 16372 26794 16552
rect 26534 16361 26587 16372
rect 26621 16361 26794 16372
rect 26534 16352 26794 16361
rect 26834 16552 27574 16572
rect 26834 16372 26854 16552
rect 26954 16372 27574 16552
rect 26834 16352 27574 16372
rect 27654 16352 27874 16572
rect 26581 16349 26627 16352
rect 26121 16312 26313 16317
rect 26379 16312 26571 16317
rect 27034 16312 27874 16352
rect 26114 16311 26574 16312
rect 26114 16277 26133 16311
rect 26301 16277 26391 16311
rect 26559 16277 26574 16311
rect 24614 16252 24754 16272
rect 24614 15812 24634 16252
rect 24734 15812 24754 16252
rect 26114 16212 26574 16277
rect 26114 16032 26134 16212
rect 26554 16032 26574 16212
rect 26114 16012 26574 16032
rect 24614 15792 24754 15812
rect 25752 15672 26764 15692
rect 25752 15612 25774 15672
rect 26734 15661 26764 15672
rect 26735 15627 26764 15661
rect 26734 15612 26764 15627
rect 25752 15596 26764 15612
rect 18814 15392 24514 15452
rect 25394 15432 26394 15452
rect 24794 15393 24994 15412
rect 24794 15392 24836 15393
rect 24942 15392 24994 15393
rect 13312 15362 13712 15382
rect 12570 15262 13582 15278
rect 22714 15270 23874 15272
rect 12570 15202 12592 15262
rect 13572 15202 13582 15262
rect 12570 15182 13582 15202
rect 22710 15252 23874 15270
rect 10832 15042 11812 15062
rect 22710 15172 22734 15252
rect 23854 15172 23874 15252
rect 22710 15152 23874 15172
rect 22710 15100 23298 15152
rect 24794 15132 24814 15392
rect 22710 14994 22838 15100
rect 23235 14994 23298 15100
rect 22710 14958 23298 14994
rect 24014 15112 24814 15132
rect 24014 14932 24034 15112
rect 24974 14932 24994 15392
rect 25394 15252 25414 15432
rect 25594 15356 26394 15432
rect 25594 15322 25896 15356
rect 26384 15322 26394 15356
rect 25594 15252 26394 15322
rect 25394 15232 26394 15252
rect 26494 15432 26894 15452
rect 26494 15420 26694 15432
rect 26494 15256 26508 15420
rect 26556 15256 26694 15420
rect 26494 15252 26694 15256
rect 26874 15252 26894 15432
rect 26494 15232 26894 15252
rect 25752 15132 26764 15148
rect 25752 15072 25774 15132
rect 26754 15072 26764 15132
rect 25752 15052 26764 15072
rect 24014 14912 24994 14932
<< via1 >>
rect 12936 38458 13356 38638
rect 25724 38576 26144 38756
rect 12716 38123 12873 38298
rect 12873 38123 12907 38298
rect 12907 38123 12936 38298
rect 12716 38118 12936 38123
rect 13356 38123 13389 38298
rect 13389 38123 13423 38298
rect 13423 38123 13576 38298
rect 13356 38118 13576 38123
rect 14556 38078 14636 38298
rect 25504 38241 25661 38416
rect 25661 38241 25695 38416
rect 25695 38241 25724 38416
rect 25504 38236 25724 38241
rect 26144 38241 26177 38416
rect 26177 38241 26211 38416
rect 26211 38241 26364 38416
rect 26144 38236 26364 38241
rect 27344 38196 27424 38416
rect 20234 38056 23444 38096
rect 7446 37938 10656 37978
rect 7446 37898 10656 37938
rect 7446 37818 10656 37898
rect 7446 37238 10606 37258
rect 7446 37198 10576 37238
rect 10576 37198 10606 37238
rect 7446 37178 10606 37198
rect 7706 36928 7748 36988
rect 7748 36928 7782 36988
rect 7782 36928 7816 36988
rect 8226 36928 8264 36988
rect 8264 36928 8298 36988
rect 8298 36928 8336 36988
rect 8736 36922 8780 36988
rect 8780 36922 8814 36988
rect 8814 36922 8846 36988
rect 8736 36878 8846 36922
rect 9256 36928 9296 36998
rect 9296 36928 9330 36998
rect 9330 36928 9366 36998
rect 9776 36922 9812 36998
rect 9812 36922 9846 36998
rect 9846 36922 9886 36998
rect 9776 36878 9886 36922
rect 10286 36928 10328 36998
rect 10328 36928 10362 36998
rect 10362 36928 10396 36998
rect 7706 36608 7748 36668
rect 7748 36608 7782 36668
rect 7782 36608 7816 36668
rect 8086 36618 8176 36778
rect 8226 36608 8264 36668
rect 8264 36608 8298 36668
rect 8298 36608 8336 36668
rect 7966 36498 8006 36558
rect 8006 36498 8040 36558
rect 8040 36498 8076 36558
rect 8486 36498 8522 36558
rect 8522 36498 8556 36558
rect 8556 36498 8596 36558
rect 8736 36608 8780 36668
rect 8780 36608 8814 36668
rect 8814 36608 8846 36668
rect 9006 36498 9038 36558
rect 9038 36498 9072 36558
rect 9072 36498 9116 36558
rect 9256 36608 9296 36668
rect 9296 36608 9330 36668
rect 9330 36608 9366 36668
rect 9516 36498 9554 36558
rect 9554 36498 9588 36558
rect 9588 36498 9626 36558
rect 9776 36608 9812 36668
rect 9812 36608 9846 36668
rect 9846 36608 9886 36668
rect 10156 36628 10236 36778
rect 10026 36498 10070 36558
rect 10070 36498 10104 36558
rect 10104 36498 10136 36558
rect 10286 36608 10328 36668
rect 10328 36608 10362 36668
rect 10362 36608 10396 36668
rect 8946 36319 9166 36368
rect 8946 36308 9010 36319
rect 9010 36308 9100 36319
rect 9100 36308 9166 36319
rect 8511 36235 8566 36248
rect 8511 36175 8522 36235
rect 8522 36175 8556 36235
rect 8556 36175 8566 36235
rect 8511 36173 8566 36175
rect 6946 36108 7366 36128
rect 6946 36018 6956 36108
rect 6956 36018 7356 36108
rect 7356 36018 7366 36108
rect 6946 36008 7366 36018
rect 9541 36235 9596 36248
rect 9541 36175 9554 36235
rect 9554 36175 9588 36235
rect 9588 36175 9596 36235
rect 9541 36173 9596 36175
rect 7506 36048 10606 36058
rect 7506 35998 7526 36048
rect 7526 35998 10576 36048
rect 10576 35998 10606 36048
rect 7506 35988 10606 35998
rect 7446 35628 10656 35678
rect 7446 35588 10656 35628
rect 7446 35518 10656 35588
rect 11596 37598 11816 37658
rect 11596 37198 11636 37598
rect 11636 37198 11756 37598
rect 11756 37198 11816 37598
rect 11596 37178 11816 37198
rect 12716 37803 12936 37818
rect 12716 37638 12873 37803
rect 12873 37638 12907 37803
rect 12907 37638 12936 37803
rect 13356 37803 13576 37818
rect 13356 37638 13389 37803
rect 13389 37638 13423 37803
rect 13423 37638 13576 37803
rect 14376 37618 14456 37838
rect 12936 37298 13356 37478
rect 12936 36998 13356 37178
rect 12716 36663 12873 36838
rect 12873 36663 12907 36838
rect 12907 36663 12936 36838
rect 12716 36658 12936 36663
rect 13356 36663 13389 36838
rect 13389 36663 13423 36838
rect 13423 36663 13576 36838
rect 13356 36658 13576 36663
rect 14556 36618 14636 36838
rect 12716 36343 12936 36358
rect 12716 36178 12873 36343
rect 12873 36178 12907 36343
rect 12907 36178 12936 36343
rect 13356 36343 13576 36358
rect 13356 36178 13389 36343
rect 13389 36178 13423 36343
rect 13423 36178 13576 36343
rect 14376 36158 14456 36378
rect 12936 35838 13356 36018
rect 12576 35467 13536 35478
rect 12576 35433 12583 35467
rect 12583 35433 12617 35467
rect 12617 35433 12675 35467
rect 12675 35433 12709 35467
rect 12709 35433 12767 35467
rect 12767 35433 12801 35467
rect 12801 35433 12859 35467
rect 12859 35433 12893 35467
rect 12893 35433 12951 35467
rect 12951 35433 12985 35467
rect 12985 35433 13043 35467
rect 13043 35433 13077 35467
rect 13077 35433 13135 35467
rect 13135 35433 13169 35467
rect 13169 35433 13227 35467
rect 13227 35433 13261 35467
rect 13261 35433 13319 35467
rect 13319 35433 13353 35467
rect 13353 35433 13411 35467
rect 13411 35433 13445 35467
rect 13445 35433 13503 35467
rect 13503 35433 13536 35467
rect 12576 35418 13536 35433
rect 20234 38016 23444 38056
rect 20234 37936 23444 38016
rect 20234 37356 23394 37376
rect 20234 37316 23364 37356
rect 23364 37316 23394 37356
rect 20234 37296 23394 37316
rect 20494 37046 20536 37106
rect 20536 37046 20570 37106
rect 20570 37046 20604 37106
rect 21014 37046 21052 37106
rect 21052 37046 21086 37106
rect 21086 37046 21124 37106
rect 21524 37040 21568 37106
rect 21568 37040 21602 37106
rect 21602 37040 21634 37106
rect 21524 36996 21634 37040
rect 22044 37046 22084 37116
rect 22084 37046 22118 37116
rect 22118 37046 22154 37116
rect 22564 37040 22600 37116
rect 22600 37040 22634 37116
rect 22634 37040 22674 37116
rect 22564 36996 22674 37040
rect 23074 37046 23116 37116
rect 23116 37046 23150 37116
rect 23150 37046 23184 37116
rect 20494 36726 20536 36786
rect 20536 36726 20570 36786
rect 20570 36726 20604 36786
rect 20874 36736 20964 36896
rect 21014 36726 21052 36786
rect 21052 36726 21086 36786
rect 21086 36726 21124 36786
rect 20754 36616 20794 36676
rect 20794 36616 20828 36676
rect 20828 36616 20864 36676
rect 21274 36616 21310 36676
rect 21310 36616 21344 36676
rect 21344 36616 21384 36676
rect 21524 36726 21568 36786
rect 21568 36726 21602 36786
rect 21602 36726 21634 36786
rect 21794 36616 21826 36676
rect 21826 36616 21860 36676
rect 21860 36616 21904 36676
rect 22044 36726 22084 36786
rect 22084 36726 22118 36786
rect 22118 36726 22154 36786
rect 22304 36616 22342 36676
rect 22342 36616 22376 36676
rect 22376 36616 22414 36676
rect 22564 36726 22600 36786
rect 22600 36726 22634 36786
rect 22634 36726 22674 36786
rect 22944 36746 23024 36896
rect 22814 36616 22858 36676
rect 22858 36616 22892 36676
rect 22892 36616 22924 36676
rect 23074 36726 23116 36786
rect 23116 36726 23150 36786
rect 23150 36726 23184 36786
rect 21734 36437 21954 36486
rect 21734 36426 21798 36437
rect 21798 36426 21888 36437
rect 21888 36426 21954 36437
rect 21299 36353 21354 36366
rect 21299 36293 21310 36353
rect 21310 36293 21344 36353
rect 21344 36293 21354 36353
rect 21299 36291 21354 36293
rect 19734 36226 20154 36246
rect 19734 36136 19744 36226
rect 19744 36136 20144 36226
rect 20144 36136 20154 36226
rect 19734 36126 20154 36136
rect 22329 36353 22384 36366
rect 22329 36293 22342 36353
rect 22342 36293 22376 36353
rect 22376 36293 22384 36353
rect 22329 36291 22384 36293
rect 20294 36166 23394 36176
rect 20294 36116 20314 36166
rect 20314 36116 23364 36166
rect 23364 36116 23394 36166
rect 20294 36106 23394 36116
rect 20234 35746 23444 35796
rect 20234 35706 23444 35746
rect 20234 35636 23444 35706
rect 24384 37716 24604 37776
rect 24384 37316 24424 37716
rect 24424 37316 24544 37716
rect 24544 37316 24604 37716
rect 24384 37296 24604 37316
rect 25504 37921 25724 37936
rect 25504 37756 25661 37921
rect 25661 37756 25695 37921
rect 25695 37756 25724 37921
rect 26144 37921 26364 37936
rect 26144 37756 26177 37921
rect 26177 37756 26211 37921
rect 26211 37756 26364 37921
rect 27164 37736 27244 37956
rect 25724 37416 26144 37596
rect 25724 37116 26144 37296
rect 25504 36781 25661 36956
rect 25661 36781 25695 36956
rect 25695 36781 25724 36956
rect 25504 36776 25724 36781
rect 26144 36781 26177 36956
rect 26177 36781 26211 36956
rect 26211 36781 26364 36956
rect 26144 36776 26364 36781
rect 27344 36736 27424 36956
rect 25504 36461 25724 36476
rect 25504 36296 25661 36461
rect 25661 36296 25695 36461
rect 25695 36296 25724 36461
rect 26144 36461 26364 36476
rect 26144 36296 26177 36461
rect 26177 36296 26211 36461
rect 26211 36296 26364 36461
rect 27164 36276 27244 36496
rect 24224 35736 24324 36176
rect 25724 35956 26144 36136
rect 25364 35585 26324 35596
rect 25364 35551 25371 35585
rect 25371 35551 25405 35585
rect 25405 35551 25463 35585
rect 25463 35551 25497 35585
rect 25497 35551 25555 35585
rect 25555 35551 25589 35585
rect 25589 35551 25647 35585
rect 25647 35551 25681 35585
rect 25681 35551 25739 35585
rect 25739 35551 25773 35585
rect 25773 35551 25831 35585
rect 25831 35551 25865 35585
rect 25865 35551 25923 35585
rect 25923 35551 25957 35585
rect 25957 35551 26015 35585
rect 26015 35551 26049 35585
rect 26049 35551 26107 35585
rect 26107 35551 26141 35585
rect 26141 35551 26199 35585
rect 26199 35551 26233 35585
rect 26233 35551 26291 35585
rect 26291 35551 26324 35585
rect 25364 35536 26324 35551
rect 12216 35058 12396 35238
rect 13496 35058 13676 35238
rect 22324 35096 23444 35176
rect 12576 34923 13556 34938
rect 12576 34889 12583 34923
rect 12583 34889 12617 34923
rect 12617 34889 12675 34923
rect 12675 34889 12709 34923
rect 12709 34889 12767 34923
rect 12767 34889 12801 34923
rect 12801 34889 12859 34923
rect 12859 34889 12893 34923
rect 12893 34889 12951 34923
rect 12951 34889 12985 34923
rect 12985 34889 13043 34923
rect 13043 34889 13077 34923
rect 13077 34889 13135 34923
rect 13135 34889 13169 34923
rect 13169 34889 13227 34923
rect 13227 34889 13261 34923
rect 13261 34889 13319 34923
rect 13319 34889 13353 34923
rect 13353 34889 13411 34923
rect 13411 34889 13445 34923
rect 13445 34889 13503 34923
rect 13503 34889 13537 34923
rect 13537 34889 13556 34923
rect 12576 34878 13556 34889
rect 24404 35036 24426 35316
rect 23624 35024 24426 35036
rect 23624 34918 23627 35024
rect 23627 34918 24024 35024
rect 24024 34920 24426 35024
rect 24426 34920 24532 35316
rect 24532 34920 24564 35316
rect 24024 34918 24564 34920
rect 23624 34856 24564 34918
rect 25004 35176 25184 35356
rect 26284 35176 26464 35356
rect 25364 35041 26344 35056
rect 25364 35007 25371 35041
rect 25371 35007 25405 35041
rect 25405 35007 25463 35041
rect 25463 35007 25497 35041
rect 25497 35007 25555 35041
rect 25555 35007 25589 35041
rect 25589 35007 25647 35041
rect 25647 35007 25681 35041
rect 25681 35007 25739 35041
rect 25739 35007 25773 35041
rect 25773 35007 25831 35041
rect 25831 35007 25865 35041
rect 25865 35007 25923 35041
rect 25923 35007 25957 35041
rect 25957 35007 26015 35041
rect 26015 35007 26049 35041
rect 26049 35007 26107 35041
rect 26107 35007 26141 35041
rect 26141 35007 26199 35041
rect 26199 35007 26233 35041
rect 26233 35007 26291 35041
rect 26291 35007 26325 35041
rect 26325 35007 26344 35041
rect 25364 34996 26344 35007
rect 12956 32532 13376 32712
rect 25688 32456 26108 32636
rect 12736 32197 12893 32372
rect 12893 32197 12927 32372
rect 12927 32197 12956 32372
rect 12736 32192 12956 32197
rect 13376 32197 13409 32372
rect 13409 32197 13443 32372
rect 13443 32197 13596 32372
rect 13376 32192 13596 32197
rect 14576 32152 14656 32372
rect 25468 32121 25625 32296
rect 25625 32121 25659 32296
rect 25659 32121 25688 32296
rect 25468 32116 25688 32121
rect 7466 32012 10676 32052
rect 7466 31972 10676 32012
rect 7466 31892 10676 31972
rect 7466 31312 10626 31332
rect 7466 31272 10596 31312
rect 10596 31272 10626 31312
rect 7466 31252 10626 31272
rect 7726 31002 7768 31062
rect 7768 31002 7802 31062
rect 7802 31002 7836 31062
rect 8246 31002 8284 31062
rect 8284 31002 8318 31062
rect 8318 31002 8356 31062
rect 8756 30996 8800 31062
rect 8800 30996 8834 31062
rect 8834 30996 8866 31062
rect 8756 30952 8866 30996
rect 9276 31002 9316 31072
rect 9316 31002 9350 31072
rect 9350 31002 9386 31072
rect 9796 30996 9832 31072
rect 9832 30996 9866 31072
rect 9866 30996 9906 31072
rect 9796 30952 9906 30996
rect 10306 31002 10348 31072
rect 10348 31002 10382 31072
rect 10382 31002 10416 31072
rect 7726 30682 7768 30742
rect 7768 30682 7802 30742
rect 7802 30682 7836 30742
rect 8106 30692 8196 30852
rect 8246 30682 8284 30742
rect 8284 30682 8318 30742
rect 8318 30682 8356 30742
rect 7986 30572 8026 30632
rect 8026 30572 8060 30632
rect 8060 30572 8096 30632
rect 8506 30572 8542 30632
rect 8542 30572 8576 30632
rect 8576 30572 8616 30632
rect 8756 30682 8800 30742
rect 8800 30682 8834 30742
rect 8834 30682 8866 30742
rect 9026 30572 9058 30632
rect 9058 30572 9092 30632
rect 9092 30572 9136 30632
rect 9276 30682 9316 30742
rect 9316 30682 9350 30742
rect 9350 30682 9386 30742
rect 9536 30572 9574 30632
rect 9574 30572 9608 30632
rect 9608 30572 9646 30632
rect 9796 30682 9832 30742
rect 9832 30682 9866 30742
rect 9866 30682 9906 30742
rect 10176 30702 10256 30852
rect 10046 30572 10090 30632
rect 10090 30572 10124 30632
rect 10124 30572 10156 30632
rect 10306 30682 10348 30742
rect 10348 30682 10382 30742
rect 10382 30682 10416 30742
rect 8966 30393 9186 30442
rect 8966 30382 9030 30393
rect 9030 30382 9120 30393
rect 9120 30382 9186 30393
rect 8531 30309 8586 30322
rect 8531 30249 8542 30309
rect 8542 30249 8576 30309
rect 8576 30249 8586 30309
rect 8531 30247 8586 30249
rect 6966 30182 7386 30202
rect 6966 30092 6976 30182
rect 6976 30092 7376 30182
rect 7376 30092 7386 30182
rect 6966 30082 7386 30092
rect 9561 30309 9616 30322
rect 9561 30249 9574 30309
rect 9574 30249 9608 30309
rect 9608 30249 9616 30309
rect 9561 30247 9616 30249
rect 7526 30122 10626 30132
rect 7526 30072 7546 30122
rect 7546 30072 10596 30122
rect 10596 30072 10626 30122
rect 7526 30062 10626 30072
rect 7466 29702 10676 29752
rect 7466 29662 10676 29702
rect 7466 29592 10676 29662
rect 26108 32121 26141 32296
rect 26141 32121 26175 32296
rect 26175 32121 26328 32296
rect 26108 32116 26328 32121
rect 27308 32076 27388 32296
rect 11616 31672 11836 31732
rect 11616 31272 11656 31672
rect 11656 31272 11776 31672
rect 11776 31272 11836 31672
rect 11616 31252 11836 31272
rect 12736 31877 12956 31892
rect 12736 31712 12893 31877
rect 12893 31712 12927 31877
rect 12927 31712 12956 31877
rect 13376 31877 13596 31892
rect 13376 31712 13409 31877
rect 13409 31712 13443 31877
rect 13443 31712 13596 31877
rect 14396 31692 14476 31912
rect 20198 31936 23408 31976
rect 12956 31372 13376 31552
rect 12956 31072 13376 31252
rect 12736 30737 12893 30912
rect 12893 30737 12927 30912
rect 12927 30737 12956 30912
rect 12736 30732 12956 30737
rect 13376 30737 13409 30912
rect 13409 30737 13443 30912
rect 13443 30737 13596 30912
rect 13376 30732 13596 30737
rect 14576 30692 14656 30912
rect 12736 30417 12956 30432
rect 12736 30252 12893 30417
rect 12893 30252 12927 30417
rect 12927 30252 12956 30417
rect 13376 30417 13596 30432
rect 13376 30252 13409 30417
rect 13409 30252 13443 30417
rect 13443 30252 13596 30417
rect 14396 30232 14476 30452
rect 11456 29692 11556 30132
rect 12956 29912 13376 30092
rect 12596 29541 13556 29552
rect 12596 29507 12603 29541
rect 12603 29507 12637 29541
rect 12637 29507 12695 29541
rect 12695 29507 12729 29541
rect 12729 29507 12787 29541
rect 12787 29507 12821 29541
rect 12821 29507 12879 29541
rect 12879 29507 12913 29541
rect 12913 29507 12971 29541
rect 12971 29507 13005 29541
rect 13005 29507 13063 29541
rect 13063 29507 13097 29541
rect 13097 29507 13155 29541
rect 13155 29507 13189 29541
rect 13189 29507 13247 29541
rect 13247 29507 13281 29541
rect 13281 29507 13339 29541
rect 13339 29507 13373 29541
rect 13373 29507 13431 29541
rect 13431 29507 13465 29541
rect 13465 29507 13523 29541
rect 13523 29507 13556 29541
rect 12596 29492 13556 29507
rect 9556 29052 10676 29132
rect 11636 28992 11658 29272
rect 10856 28980 11658 28992
rect 10856 28874 10859 28980
rect 10859 28874 11256 28980
rect 11256 28876 11658 28980
rect 11658 28876 11764 29272
rect 11764 28876 11796 29272
rect 11256 28874 11796 28876
rect 10856 28812 11796 28874
rect 12236 29132 12416 29312
rect 13516 29132 13696 29312
rect 20198 31896 23408 31936
rect 20198 31816 23408 31896
rect 20198 31236 23358 31256
rect 20198 31196 23328 31236
rect 23328 31196 23358 31236
rect 20198 31176 23358 31196
rect 20458 30926 20500 30986
rect 20500 30926 20534 30986
rect 20534 30926 20568 30986
rect 20978 30926 21016 30986
rect 21016 30926 21050 30986
rect 21050 30926 21088 30986
rect 21488 30920 21532 30986
rect 21532 30920 21566 30986
rect 21566 30920 21598 30986
rect 21488 30876 21598 30920
rect 22008 30926 22048 30996
rect 22048 30926 22082 30996
rect 22082 30926 22118 30996
rect 22528 30920 22564 30996
rect 22564 30920 22598 30996
rect 22598 30920 22638 30996
rect 22528 30876 22638 30920
rect 23038 30926 23080 30996
rect 23080 30926 23114 30996
rect 23114 30926 23148 30996
rect 20458 30606 20500 30666
rect 20500 30606 20534 30666
rect 20534 30606 20568 30666
rect 20838 30616 20928 30776
rect 20978 30606 21016 30666
rect 21016 30606 21050 30666
rect 21050 30606 21088 30666
rect 20718 30496 20758 30556
rect 20758 30496 20792 30556
rect 20792 30496 20828 30556
rect 21238 30496 21274 30556
rect 21274 30496 21308 30556
rect 21308 30496 21348 30556
rect 21488 30606 21532 30666
rect 21532 30606 21566 30666
rect 21566 30606 21598 30666
rect 21758 30496 21790 30556
rect 21790 30496 21824 30556
rect 21824 30496 21868 30556
rect 22008 30606 22048 30666
rect 22048 30606 22082 30666
rect 22082 30606 22118 30666
rect 22268 30496 22306 30556
rect 22306 30496 22340 30556
rect 22340 30496 22378 30556
rect 22528 30606 22564 30666
rect 22564 30606 22598 30666
rect 22598 30606 22638 30666
rect 22908 30626 22988 30776
rect 22778 30496 22822 30556
rect 22822 30496 22856 30556
rect 22856 30496 22888 30556
rect 23038 30606 23080 30666
rect 23080 30606 23114 30666
rect 23114 30606 23148 30666
rect 21698 30317 21918 30366
rect 21698 30306 21762 30317
rect 21762 30306 21852 30317
rect 21852 30306 21918 30317
rect 21263 30233 21318 30246
rect 21263 30173 21274 30233
rect 21274 30173 21308 30233
rect 21308 30173 21318 30233
rect 21263 30171 21318 30173
rect 19698 30106 20118 30126
rect 19698 30016 19708 30106
rect 19708 30016 20108 30106
rect 20108 30016 20118 30106
rect 19698 30006 20118 30016
rect 22293 30233 22348 30246
rect 22293 30173 22306 30233
rect 22306 30173 22340 30233
rect 22340 30173 22348 30233
rect 22293 30171 22348 30173
rect 20258 30046 23358 30056
rect 20258 29996 20278 30046
rect 20278 29996 23328 30046
rect 23328 29996 23358 30046
rect 20258 29986 23358 29996
rect 20198 29626 23408 29676
rect 20198 29586 23408 29626
rect 20198 29516 23408 29586
rect 24348 31596 24568 31656
rect 24348 31196 24388 31596
rect 24388 31196 24508 31596
rect 24508 31196 24568 31596
rect 24348 31176 24568 31196
rect 25468 31801 25688 31816
rect 25468 31636 25625 31801
rect 25625 31636 25659 31801
rect 25659 31636 25688 31801
rect 26108 31801 26328 31816
rect 26108 31636 26141 31801
rect 26141 31636 26175 31801
rect 26175 31636 26328 31801
rect 27128 31616 27208 31836
rect 25688 31296 26108 31476
rect 25688 30996 26108 31176
rect 25468 30661 25625 30836
rect 25625 30661 25659 30836
rect 25659 30661 25688 30836
rect 25468 30656 25688 30661
rect 26108 30661 26141 30836
rect 26141 30661 26175 30836
rect 26175 30661 26328 30836
rect 26108 30656 26328 30661
rect 27308 30616 27388 30836
rect 25468 30341 25688 30356
rect 25468 30176 25625 30341
rect 25625 30176 25659 30341
rect 25659 30176 25688 30341
rect 26108 30341 26328 30356
rect 26108 30176 26141 30341
rect 26141 30176 26175 30341
rect 26175 30176 26328 30341
rect 27128 30156 27208 30376
rect 24188 29616 24288 30056
rect 25688 29836 26108 30016
rect 25328 29465 26288 29476
rect 25328 29431 25335 29465
rect 25335 29431 25369 29465
rect 25369 29431 25427 29465
rect 25427 29431 25461 29465
rect 25461 29431 25519 29465
rect 25519 29431 25553 29465
rect 25553 29431 25611 29465
rect 25611 29431 25645 29465
rect 25645 29431 25703 29465
rect 25703 29431 25737 29465
rect 25737 29431 25795 29465
rect 25795 29431 25829 29465
rect 25829 29431 25887 29465
rect 25887 29431 25921 29465
rect 25921 29431 25979 29465
rect 25979 29431 26013 29465
rect 26013 29431 26071 29465
rect 26071 29431 26105 29465
rect 26105 29431 26163 29465
rect 26163 29431 26197 29465
rect 26197 29431 26255 29465
rect 26255 29431 26288 29465
rect 25328 29416 26288 29431
rect 12596 28997 13576 29012
rect 12596 28963 12603 28997
rect 12603 28963 12637 28997
rect 12637 28963 12695 28997
rect 12695 28963 12729 28997
rect 12729 28963 12787 28997
rect 12787 28963 12821 28997
rect 12821 28963 12879 28997
rect 12879 28963 12913 28997
rect 12913 28963 12971 28997
rect 12971 28963 13005 28997
rect 13005 28963 13063 28997
rect 13063 28963 13097 28997
rect 13097 28963 13155 28997
rect 13155 28963 13189 28997
rect 13189 28963 13247 28997
rect 13247 28963 13281 28997
rect 13281 28963 13339 28997
rect 13339 28963 13373 28997
rect 13373 28963 13431 28997
rect 13431 28963 13465 28997
rect 13465 28963 13523 28997
rect 13523 28963 13557 28997
rect 13557 28963 13576 28997
rect 12596 28952 13576 28963
rect 22288 28976 23408 29056
rect 24368 28916 24390 29196
rect 23588 28904 24390 28916
rect 23588 28798 23591 28904
rect 23591 28798 23988 28904
rect 23988 28800 24390 28904
rect 24390 28800 24496 29196
rect 24496 28800 24528 29196
rect 23988 28798 24528 28800
rect 23588 28736 24528 28798
rect 24968 29056 25148 29236
rect 26248 29056 26428 29236
rect 25328 28921 26308 28936
rect 25328 28887 25335 28921
rect 25335 28887 25369 28921
rect 25369 28887 25427 28921
rect 25427 28887 25461 28921
rect 25461 28887 25519 28921
rect 25519 28887 25553 28921
rect 25553 28887 25611 28921
rect 25611 28887 25645 28921
rect 25645 28887 25703 28921
rect 25703 28887 25737 28921
rect 25737 28887 25795 28921
rect 25795 28887 25829 28921
rect 25829 28887 25887 28921
rect 25887 28887 25921 28921
rect 25921 28887 25979 28921
rect 25979 28887 26013 28921
rect 26013 28887 26071 28921
rect 26071 28887 26105 28921
rect 26105 28887 26163 28921
rect 26163 28887 26197 28921
rect 26197 28887 26255 28921
rect 26255 28887 26289 28921
rect 26289 28887 26308 28921
rect 25328 28876 26308 28887
rect 13076 25828 13496 26008
rect 12856 25493 13013 25668
rect 13013 25493 13047 25668
rect 13047 25493 13076 25668
rect 12856 25488 13076 25493
rect 13496 25493 13529 25668
rect 13529 25493 13563 25668
rect 13563 25493 13716 25668
rect 13496 25488 13716 25493
rect 14696 25448 14776 25668
rect 25784 25698 26204 25878
rect 7586 25308 10796 25348
rect 7586 25268 10796 25308
rect 7586 25188 10796 25268
rect 7586 24608 10746 24628
rect 7586 24568 10716 24608
rect 10716 24568 10746 24608
rect 7586 24548 10746 24568
rect 7846 24298 7888 24358
rect 7888 24298 7922 24358
rect 7922 24298 7956 24358
rect 8366 24298 8404 24358
rect 8404 24298 8438 24358
rect 8438 24298 8476 24358
rect 8876 24292 8920 24358
rect 8920 24292 8954 24358
rect 8954 24292 8986 24358
rect 8876 24248 8986 24292
rect 9396 24298 9436 24368
rect 9436 24298 9470 24368
rect 9470 24298 9506 24368
rect 9916 24292 9952 24368
rect 9952 24292 9986 24368
rect 9986 24292 10026 24368
rect 9916 24248 10026 24292
rect 10426 24298 10468 24368
rect 10468 24298 10502 24368
rect 10502 24298 10536 24368
rect 7846 23978 7888 24038
rect 7888 23978 7922 24038
rect 7922 23978 7956 24038
rect 8226 23988 8316 24148
rect 8366 23978 8404 24038
rect 8404 23978 8438 24038
rect 8438 23978 8476 24038
rect 8106 23868 8146 23928
rect 8146 23868 8180 23928
rect 8180 23868 8216 23928
rect 8626 23868 8662 23928
rect 8662 23868 8696 23928
rect 8696 23868 8736 23928
rect 8876 23978 8920 24038
rect 8920 23978 8954 24038
rect 8954 23978 8986 24038
rect 9146 23868 9178 23928
rect 9178 23868 9212 23928
rect 9212 23868 9256 23928
rect 9396 23978 9436 24038
rect 9436 23978 9470 24038
rect 9470 23978 9506 24038
rect 9656 23868 9694 23928
rect 9694 23868 9728 23928
rect 9728 23868 9766 23928
rect 9916 23978 9952 24038
rect 9952 23978 9986 24038
rect 9986 23978 10026 24038
rect 10296 23998 10376 24148
rect 10166 23868 10210 23928
rect 10210 23868 10244 23928
rect 10244 23868 10276 23928
rect 10426 23978 10468 24038
rect 10468 23978 10502 24038
rect 10502 23978 10536 24038
rect 9086 23689 9306 23738
rect 9086 23678 9150 23689
rect 9150 23678 9240 23689
rect 9240 23678 9306 23689
rect 8651 23605 8706 23618
rect 8651 23545 8662 23605
rect 8662 23545 8696 23605
rect 8696 23545 8706 23605
rect 8651 23543 8706 23545
rect 7086 23478 7506 23498
rect 7086 23388 7096 23478
rect 7096 23388 7496 23478
rect 7496 23388 7506 23478
rect 7086 23378 7506 23388
rect 9681 23605 9736 23618
rect 9681 23545 9694 23605
rect 9694 23545 9728 23605
rect 9728 23545 9736 23605
rect 9681 23543 9736 23545
rect 7646 23418 10746 23428
rect 7646 23368 7666 23418
rect 7666 23368 10716 23418
rect 10716 23368 10746 23418
rect 7646 23358 10746 23368
rect 7586 22998 10796 23048
rect 7586 22958 10796 22998
rect 7586 22888 10796 22958
rect 25564 25363 25721 25538
rect 25721 25363 25755 25538
rect 25755 25363 25784 25538
rect 25564 25358 25784 25363
rect 26204 25363 26237 25538
rect 26237 25363 26271 25538
rect 26271 25363 26424 25538
rect 26204 25358 26424 25363
rect 27404 25318 27484 25538
rect 11736 24968 11956 25028
rect 11736 24568 11776 24968
rect 11776 24568 11896 24968
rect 11896 24568 11956 24968
rect 11736 24548 11956 24568
rect 12856 25173 13076 25188
rect 12856 25008 13013 25173
rect 13013 25008 13047 25173
rect 13047 25008 13076 25173
rect 13496 25173 13716 25188
rect 13496 25008 13529 25173
rect 13529 25008 13563 25173
rect 13563 25008 13716 25173
rect 14516 24988 14596 25208
rect 20294 25178 23504 25218
rect 13076 24668 13496 24848
rect 13076 24368 13496 24548
rect 12856 24033 13013 24208
rect 13013 24033 13047 24208
rect 13047 24033 13076 24208
rect 12856 24028 13076 24033
rect 13496 24033 13529 24208
rect 13529 24033 13563 24208
rect 13563 24033 13716 24208
rect 13496 24028 13716 24033
rect 14696 23988 14776 24208
rect 12856 23713 13076 23728
rect 12856 23548 13013 23713
rect 13013 23548 13047 23713
rect 13047 23548 13076 23713
rect 13496 23713 13716 23728
rect 13496 23548 13529 23713
rect 13529 23548 13563 23713
rect 13563 23548 13716 23713
rect 14516 23528 14596 23748
rect 11576 22988 11676 23428
rect 13076 23208 13496 23388
rect 12716 22837 13676 22848
rect 12716 22803 12723 22837
rect 12723 22803 12757 22837
rect 12757 22803 12815 22837
rect 12815 22803 12849 22837
rect 12849 22803 12907 22837
rect 12907 22803 12941 22837
rect 12941 22803 12999 22837
rect 12999 22803 13033 22837
rect 13033 22803 13091 22837
rect 13091 22803 13125 22837
rect 13125 22803 13183 22837
rect 13183 22803 13217 22837
rect 13217 22803 13275 22837
rect 13275 22803 13309 22837
rect 13309 22803 13367 22837
rect 13367 22803 13401 22837
rect 13401 22803 13459 22837
rect 13459 22803 13493 22837
rect 13493 22803 13551 22837
rect 13551 22803 13585 22837
rect 13585 22803 13643 22837
rect 13643 22803 13676 22837
rect 12716 22788 13676 22803
rect 9676 22348 10796 22428
rect 11756 22288 11778 22568
rect 10976 22276 11778 22288
rect 10976 22170 10979 22276
rect 10979 22170 11376 22276
rect 11376 22172 11778 22276
rect 11778 22172 11884 22568
rect 11884 22172 11916 22568
rect 11376 22170 11916 22172
rect 10976 22108 11916 22170
rect 12356 22428 12536 22608
rect 13636 22428 13816 22608
rect 20294 25138 23504 25178
rect 20294 25058 23504 25138
rect 20294 24478 23454 24498
rect 20294 24438 23424 24478
rect 23424 24438 23454 24478
rect 20294 24418 23454 24438
rect 20554 24168 20596 24228
rect 20596 24168 20630 24228
rect 20630 24168 20664 24228
rect 21074 24168 21112 24228
rect 21112 24168 21146 24228
rect 21146 24168 21184 24228
rect 21584 24162 21628 24228
rect 21628 24162 21662 24228
rect 21662 24162 21694 24228
rect 21584 24118 21694 24162
rect 22104 24168 22144 24238
rect 22144 24168 22178 24238
rect 22178 24168 22214 24238
rect 22624 24162 22660 24238
rect 22660 24162 22694 24238
rect 22694 24162 22734 24238
rect 22624 24118 22734 24162
rect 23134 24168 23176 24238
rect 23176 24168 23210 24238
rect 23210 24168 23244 24238
rect 20554 23848 20596 23908
rect 20596 23848 20630 23908
rect 20630 23848 20664 23908
rect 20934 23858 21024 24018
rect 21074 23848 21112 23908
rect 21112 23848 21146 23908
rect 21146 23848 21184 23908
rect 20814 23738 20854 23798
rect 20854 23738 20888 23798
rect 20888 23738 20924 23798
rect 21334 23738 21370 23798
rect 21370 23738 21404 23798
rect 21404 23738 21444 23798
rect 21584 23848 21628 23908
rect 21628 23848 21662 23908
rect 21662 23848 21694 23908
rect 21854 23738 21886 23798
rect 21886 23738 21920 23798
rect 21920 23738 21964 23798
rect 22104 23848 22144 23908
rect 22144 23848 22178 23908
rect 22178 23848 22214 23908
rect 22364 23738 22402 23798
rect 22402 23738 22436 23798
rect 22436 23738 22474 23798
rect 22624 23848 22660 23908
rect 22660 23848 22694 23908
rect 22694 23848 22734 23908
rect 23004 23868 23084 24018
rect 22874 23738 22918 23798
rect 22918 23738 22952 23798
rect 22952 23738 22984 23798
rect 23134 23848 23176 23908
rect 23176 23848 23210 23908
rect 23210 23848 23244 23908
rect 21794 23559 22014 23608
rect 21794 23548 21858 23559
rect 21858 23548 21948 23559
rect 21948 23548 22014 23559
rect 21359 23475 21414 23488
rect 21359 23415 21370 23475
rect 21370 23415 21404 23475
rect 21404 23415 21414 23475
rect 21359 23413 21414 23415
rect 19794 23348 20214 23368
rect 19794 23258 19804 23348
rect 19804 23258 20204 23348
rect 20204 23258 20214 23348
rect 19794 23248 20214 23258
rect 22389 23475 22444 23488
rect 22389 23415 22402 23475
rect 22402 23415 22436 23475
rect 22436 23415 22444 23475
rect 22389 23413 22444 23415
rect 20354 23288 23454 23298
rect 20354 23238 20374 23288
rect 20374 23238 23424 23288
rect 23424 23238 23454 23288
rect 20354 23228 23454 23238
rect 20294 22868 23504 22918
rect 20294 22828 23504 22868
rect 20294 22758 23504 22828
rect 24444 24838 24664 24898
rect 24444 24438 24484 24838
rect 24484 24438 24604 24838
rect 24604 24438 24664 24838
rect 24444 24418 24664 24438
rect 25564 25043 25784 25058
rect 25564 24878 25721 25043
rect 25721 24878 25755 25043
rect 25755 24878 25784 25043
rect 26204 25043 26424 25058
rect 26204 24878 26237 25043
rect 26237 24878 26271 25043
rect 26271 24878 26424 25043
rect 27224 24858 27304 25078
rect 25784 24538 26204 24718
rect 25784 24238 26204 24418
rect 25564 23903 25721 24078
rect 25721 23903 25755 24078
rect 25755 23903 25784 24078
rect 25564 23898 25784 23903
rect 26204 23903 26237 24078
rect 26237 23903 26271 24078
rect 26271 23903 26424 24078
rect 26204 23898 26424 23903
rect 27404 23858 27484 24078
rect 25564 23583 25784 23598
rect 25564 23418 25721 23583
rect 25721 23418 25755 23583
rect 25755 23418 25784 23583
rect 26204 23583 26424 23598
rect 26204 23418 26237 23583
rect 26237 23418 26271 23583
rect 26271 23418 26424 23583
rect 27224 23398 27304 23618
rect 24284 22858 24384 23298
rect 25784 23078 26204 23258
rect 25424 22707 26384 22718
rect 25424 22673 25431 22707
rect 25431 22673 25465 22707
rect 25465 22673 25523 22707
rect 25523 22673 25557 22707
rect 25557 22673 25615 22707
rect 25615 22673 25649 22707
rect 25649 22673 25707 22707
rect 25707 22673 25741 22707
rect 25741 22673 25799 22707
rect 25799 22673 25833 22707
rect 25833 22673 25891 22707
rect 25891 22673 25925 22707
rect 25925 22673 25983 22707
rect 25983 22673 26017 22707
rect 26017 22673 26075 22707
rect 26075 22673 26109 22707
rect 26109 22673 26167 22707
rect 26167 22673 26201 22707
rect 26201 22673 26259 22707
rect 26259 22673 26293 22707
rect 26293 22673 26351 22707
rect 26351 22673 26384 22707
rect 25424 22658 26384 22673
rect 12716 22293 13696 22308
rect 12716 22259 12723 22293
rect 12723 22259 12757 22293
rect 12757 22259 12815 22293
rect 12815 22259 12849 22293
rect 12849 22259 12907 22293
rect 12907 22259 12941 22293
rect 12941 22259 12999 22293
rect 12999 22259 13033 22293
rect 13033 22259 13091 22293
rect 13091 22259 13125 22293
rect 13125 22259 13183 22293
rect 13183 22259 13217 22293
rect 13217 22259 13275 22293
rect 13275 22259 13309 22293
rect 13309 22259 13367 22293
rect 13367 22259 13401 22293
rect 13401 22259 13459 22293
rect 13459 22259 13493 22293
rect 13493 22259 13551 22293
rect 13551 22259 13585 22293
rect 13585 22259 13643 22293
rect 13643 22259 13677 22293
rect 13677 22259 13696 22293
rect 12716 22248 13696 22259
rect 22384 22218 23504 22298
rect 24464 22158 24486 22438
rect 23684 22146 24486 22158
rect 23684 22040 23687 22146
rect 23687 22040 24084 22146
rect 24084 22042 24486 22146
rect 24486 22042 24592 22438
rect 24592 22042 24624 22438
rect 24084 22040 24624 22042
rect 23684 21978 24624 22040
rect 25064 22298 25244 22478
rect 26344 22298 26524 22478
rect 25424 22163 26404 22178
rect 25424 22129 25431 22163
rect 25431 22129 25465 22163
rect 25465 22129 25523 22163
rect 25523 22129 25557 22163
rect 25557 22129 25615 22163
rect 25615 22129 25649 22163
rect 25649 22129 25707 22163
rect 25707 22129 25741 22163
rect 25741 22129 25799 22163
rect 25799 22129 25833 22163
rect 25833 22129 25891 22163
rect 25891 22129 25925 22163
rect 25925 22129 25983 22163
rect 25983 22129 26017 22163
rect 26017 22129 26075 22163
rect 26075 22129 26109 22163
rect 26109 22129 26167 22163
rect 26167 22129 26201 22163
rect 26201 22129 26259 22163
rect 26259 22129 26293 22163
rect 26293 22129 26351 22163
rect 26351 22129 26385 22163
rect 26385 22129 26404 22163
rect 25424 22118 26404 22129
rect 12952 18782 13372 18962
rect 12732 18447 12889 18622
rect 12889 18447 12923 18622
rect 12923 18447 12952 18622
rect 12732 18442 12952 18447
rect 13372 18447 13405 18622
rect 13405 18447 13439 18622
rect 13439 18447 13592 18622
rect 13372 18442 13592 18447
rect 14572 18402 14652 18622
rect 26134 18652 26554 18832
rect 7462 18262 10672 18302
rect 7462 18222 10672 18262
rect 7462 18142 10672 18222
rect 7462 17562 10622 17582
rect 7462 17522 10592 17562
rect 10592 17522 10622 17562
rect 7462 17502 10622 17522
rect 7722 17252 7764 17312
rect 7764 17252 7798 17312
rect 7798 17252 7832 17312
rect 8242 17252 8280 17312
rect 8280 17252 8314 17312
rect 8314 17252 8352 17312
rect 8752 17246 8796 17312
rect 8796 17246 8830 17312
rect 8830 17246 8862 17312
rect 8752 17202 8862 17246
rect 9272 17252 9312 17322
rect 9312 17252 9346 17322
rect 9346 17252 9382 17322
rect 9792 17246 9828 17322
rect 9828 17246 9862 17322
rect 9862 17246 9902 17322
rect 9792 17202 9902 17246
rect 10302 17252 10344 17322
rect 10344 17252 10378 17322
rect 10378 17252 10412 17322
rect 7722 16932 7764 16992
rect 7764 16932 7798 16992
rect 7798 16932 7832 16992
rect 8102 16942 8192 17102
rect 8242 16932 8280 16992
rect 8280 16932 8314 16992
rect 8314 16932 8352 16992
rect 7982 16822 8022 16882
rect 8022 16822 8056 16882
rect 8056 16822 8092 16882
rect 8502 16822 8538 16882
rect 8538 16822 8572 16882
rect 8572 16822 8612 16882
rect 8752 16932 8796 16992
rect 8796 16932 8830 16992
rect 8830 16932 8862 16992
rect 9022 16822 9054 16882
rect 9054 16822 9088 16882
rect 9088 16822 9132 16882
rect 9272 16932 9312 16992
rect 9312 16932 9346 16992
rect 9346 16932 9382 16992
rect 9532 16822 9570 16882
rect 9570 16822 9604 16882
rect 9604 16822 9642 16882
rect 9792 16932 9828 16992
rect 9828 16932 9862 16992
rect 9862 16932 9902 16992
rect 10172 16952 10252 17102
rect 10042 16822 10086 16882
rect 10086 16822 10120 16882
rect 10120 16822 10152 16882
rect 10302 16932 10344 16992
rect 10344 16932 10378 16992
rect 10378 16932 10412 16992
rect 8962 16643 9182 16692
rect 8962 16632 9026 16643
rect 9026 16632 9116 16643
rect 9116 16632 9182 16643
rect 8527 16559 8582 16572
rect 8527 16499 8538 16559
rect 8538 16499 8572 16559
rect 8572 16499 8582 16559
rect 8527 16497 8582 16499
rect 6962 16432 7382 16452
rect 6962 16342 6972 16432
rect 6972 16342 7372 16432
rect 7372 16342 7382 16432
rect 6962 16332 7382 16342
rect 9557 16559 9612 16572
rect 9557 16499 9570 16559
rect 9570 16499 9604 16559
rect 9604 16499 9612 16559
rect 9557 16497 9612 16499
rect 7522 16372 10622 16382
rect 7522 16322 7542 16372
rect 7542 16322 10592 16372
rect 10592 16322 10622 16372
rect 7522 16312 10622 16322
rect 7462 15952 10672 16002
rect 7462 15912 10672 15952
rect 7462 15842 10672 15912
rect 25914 18317 26071 18492
rect 26071 18317 26105 18492
rect 26105 18317 26134 18492
rect 25914 18312 26134 18317
rect 26554 18317 26587 18492
rect 26587 18317 26621 18492
rect 26621 18317 26774 18492
rect 26554 18312 26774 18317
rect 27754 18272 27834 18492
rect 11612 17922 11832 17982
rect 11612 17522 11652 17922
rect 11652 17522 11772 17922
rect 11772 17522 11832 17922
rect 11612 17502 11832 17522
rect 12732 18127 12952 18142
rect 12732 17962 12889 18127
rect 12889 17962 12923 18127
rect 12923 17962 12952 18127
rect 13372 18127 13592 18142
rect 13372 17962 13405 18127
rect 13405 17962 13439 18127
rect 13439 17962 13592 18127
rect 14392 17942 14472 18162
rect 20644 18132 23854 18172
rect 12952 17622 13372 17802
rect 12952 17322 13372 17502
rect 12732 16987 12889 17162
rect 12889 16987 12923 17162
rect 12923 16987 12952 17162
rect 12732 16982 12952 16987
rect 13372 16987 13405 17162
rect 13405 16987 13439 17162
rect 13439 16987 13592 17162
rect 13372 16982 13592 16987
rect 14572 16942 14652 17162
rect 12732 16667 12952 16682
rect 12732 16502 12889 16667
rect 12889 16502 12923 16667
rect 12923 16502 12952 16667
rect 13372 16667 13592 16682
rect 13372 16502 13405 16667
rect 13405 16502 13439 16667
rect 13439 16502 13592 16667
rect 14392 16482 14472 16702
rect 11452 15942 11552 16382
rect 12952 16162 13372 16342
rect 12592 15791 13552 15802
rect 12592 15757 12599 15791
rect 12599 15757 12633 15791
rect 12633 15757 12691 15791
rect 12691 15757 12725 15791
rect 12725 15757 12783 15791
rect 12783 15757 12817 15791
rect 12817 15757 12875 15791
rect 12875 15757 12909 15791
rect 12909 15757 12967 15791
rect 12967 15757 13001 15791
rect 13001 15757 13059 15791
rect 13059 15757 13093 15791
rect 13093 15757 13151 15791
rect 13151 15757 13185 15791
rect 13185 15757 13243 15791
rect 13243 15757 13277 15791
rect 13277 15757 13335 15791
rect 13335 15757 13369 15791
rect 13369 15757 13427 15791
rect 13427 15757 13461 15791
rect 13461 15757 13519 15791
rect 13519 15757 13552 15791
rect 12592 15742 13552 15757
rect 9552 15302 10672 15382
rect 11632 15242 11654 15522
rect 10852 15230 11654 15242
rect 10852 15124 10855 15230
rect 10855 15124 11252 15230
rect 11252 15126 11654 15230
rect 11654 15126 11760 15522
rect 11760 15126 11792 15522
rect 11252 15124 11792 15126
rect 10852 15062 11792 15124
rect 12232 15382 12412 15562
rect 13512 15382 13692 15562
rect 20644 18092 23854 18132
rect 20644 18012 23854 18092
rect 20644 17432 23804 17452
rect 20644 17392 23774 17432
rect 23774 17392 23804 17432
rect 20644 17372 23804 17392
rect 20904 17122 20946 17182
rect 20946 17122 20980 17182
rect 20980 17122 21014 17182
rect 21424 17122 21462 17182
rect 21462 17122 21496 17182
rect 21496 17122 21534 17182
rect 21934 17116 21978 17182
rect 21978 17116 22012 17182
rect 22012 17116 22044 17182
rect 21934 17072 22044 17116
rect 22454 17122 22494 17192
rect 22494 17122 22528 17192
rect 22528 17122 22564 17192
rect 22974 17116 23010 17192
rect 23010 17116 23044 17192
rect 23044 17116 23084 17192
rect 22974 17072 23084 17116
rect 23484 17122 23526 17192
rect 23526 17122 23560 17192
rect 23560 17122 23594 17192
rect 20904 16802 20946 16862
rect 20946 16802 20980 16862
rect 20980 16802 21014 16862
rect 21284 16812 21374 16972
rect 21424 16802 21462 16862
rect 21462 16802 21496 16862
rect 21496 16802 21534 16862
rect 21164 16692 21204 16752
rect 21204 16692 21238 16752
rect 21238 16692 21274 16752
rect 21684 16692 21720 16752
rect 21720 16692 21754 16752
rect 21754 16692 21794 16752
rect 21934 16802 21978 16862
rect 21978 16802 22012 16862
rect 22012 16802 22044 16862
rect 22204 16692 22236 16752
rect 22236 16692 22270 16752
rect 22270 16692 22314 16752
rect 22454 16802 22494 16862
rect 22494 16802 22528 16862
rect 22528 16802 22564 16862
rect 22714 16692 22752 16752
rect 22752 16692 22786 16752
rect 22786 16692 22824 16752
rect 22974 16802 23010 16862
rect 23010 16802 23044 16862
rect 23044 16802 23084 16862
rect 23354 16822 23434 16972
rect 23224 16692 23268 16752
rect 23268 16692 23302 16752
rect 23302 16692 23334 16752
rect 23484 16802 23526 16862
rect 23526 16802 23560 16862
rect 23560 16802 23594 16862
rect 22144 16513 22364 16562
rect 22144 16502 22208 16513
rect 22208 16502 22298 16513
rect 22298 16502 22364 16513
rect 21709 16429 21764 16442
rect 21709 16369 21720 16429
rect 21720 16369 21754 16429
rect 21754 16369 21764 16429
rect 21709 16367 21764 16369
rect 20144 16302 20564 16322
rect 20144 16212 20154 16302
rect 20154 16212 20554 16302
rect 20554 16212 20564 16302
rect 20144 16202 20564 16212
rect 22739 16429 22794 16442
rect 22739 16369 22752 16429
rect 22752 16369 22786 16429
rect 22786 16369 22794 16429
rect 22739 16367 22794 16369
rect 20704 16242 23804 16252
rect 20704 16192 20724 16242
rect 20724 16192 23774 16242
rect 23774 16192 23804 16242
rect 20704 16182 23804 16192
rect 20644 15822 23854 15872
rect 20644 15782 23854 15822
rect 20644 15712 23854 15782
rect 24794 17792 25014 17852
rect 24794 17392 24834 17792
rect 24834 17392 24954 17792
rect 24954 17392 25014 17792
rect 24794 17372 25014 17392
rect 25914 17997 26134 18012
rect 25914 17832 26071 17997
rect 26071 17832 26105 17997
rect 26105 17832 26134 17997
rect 26554 17997 26774 18012
rect 26554 17832 26587 17997
rect 26587 17832 26621 17997
rect 26621 17832 26774 17997
rect 27574 17812 27654 18032
rect 26134 17492 26554 17672
rect 26134 17192 26554 17372
rect 25914 16857 26071 17032
rect 26071 16857 26105 17032
rect 26105 16857 26134 17032
rect 25914 16852 26134 16857
rect 26554 16857 26587 17032
rect 26587 16857 26621 17032
rect 26621 16857 26774 17032
rect 26554 16852 26774 16857
rect 27754 16812 27834 17032
rect 25914 16537 26134 16552
rect 25914 16372 26071 16537
rect 26071 16372 26105 16537
rect 26105 16372 26134 16537
rect 26554 16537 26774 16552
rect 26554 16372 26587 16537
rect 26587 16372 26621 16537
rect 26621 16372 26774 16537
rect 27574 16352 27654 16572
rect 24634 15812 24734 16252
rect 26134 16032 26554 16212
rect 25774 15661 26734 15672
rect 25774 15627 25781 15661
rect 25781 15627 25815 15661
rect 25815 15627 25873 15661
rect 25873 15627 25907 15661
rect 25907 15627 25965 15661
rect 25965 15627 25999 15661
rect 25999 15627 26057 15661
rect 26057 15627 26091 15661
rect 26091 15627 26149 15661
rect 26149 15627 26183 15661
rect 26183 15627 26241 15661
rect 26241 15627 26275 15661
rect 26275 15627 26333 15661
rect 26333 15627 26367 15661
rect 26367 15627 26425 15661
rect 26425 15627 26459 15661
rect 26459 15627 26517 15661
rect 26517 15627 26551 15661
rect 26551 15627 26609 15661
rect 26609 15627 26643 15661
rect 26643 15627 26701 15661
rect 26701 15627 26734 15661
rect 25774 15612 26734 15627
rect 12592 15247 13572 15262
rect 12592 15213 12599 15247
rect 12599 15213 12633 15247
rect 12633 15213 12691 15247
rect 12691 15213 12725 15247
rect 12725 15213 12783 15247
rect 12783 15213 12817 15247
rect 12817 15213 12875 15247
rect 12875 15213 12909 15247
rect 12909 15213 12967 15247
rect 12967 15213 13001 15247
rect 13001 15213 13059 15247
rect 13059 15213 13093 15247
rect 13093 15213 13151 15247
rect 13151 15213 13185 15247
rect 13185 15213 13243 15247
rect 13243 15213 13277 15247
rect 13277 15213 13335 15247
rect 13335 15213 13369 15247
rect 13369 15213 13427 15247
rect 13427 15213 13461 15247
rect 13461 15213 13519 15247
rect 13519 15213 13553 15247
rect 13553 15213 13572 15247
rect 12592 15202 13572 15213
rect 22734 15172 23854 15252
rect 24814 15112 24836 15392
rect 24034 15100 24836 15112
rect 24034 14994 24037 15100
rect 24037 14994 24434 15100
rect 24434 14996 24836 15100
rect 24836 14996 24942 15392
rect 24942 14996 24974 15392
rect 24434 14994 24974 14996
rect 24034 14932 24974 14994
rect 25414 15252 25594 15432
rect 26694 15252 26874 15432
rect 25774 15117 26754 15132
rect 25774 15083 25781 15117
rect 25781 15083 25815 15117
rect 25815 15083 25873 15117
rect 25873 15083 25907 15117
rect 25907 15083 25965 15117
rect 25965 15083 25999 15117
rect 25999 15083 26057 15117
rect 26057 15083 26091 15117
rect 26091 15083 26149 15117
rect 26149 15083 26183 15117
rect 26183 15083 26241 15117
rect 26241 15083 26275 15117
rect 26275 15083 26333 15117
rect 26333 15083 26367 15117
rect 26367 15083 26425 15117
rect 26425 15083 26459 15117
rect 26459 15083 26517 15117
rect 26517 15083 26551 15117
rect 26551 15083 26609 15117
rect 26609 15083 26643 15117
rect 26643 15083 26701 15117
rect 26701 15083 26735 15117
rect 26735 15083 26754 15117
rect 25774 15072 26754 15083
<< metal2 >>
rect 14960 44600 15140 44620
rect 14960 44480 14980 44600
rect 15120 44480 15140 44600
rect 14960 44460 15140 44480
rect 15000 39944 15100 44460
rect 17380 44400 17600 44420
rect 17380 44280 17400 44400
rect 17580 44280 17600 44400
rect 17380 44260 17600 44280
rect 15380 44200 15600 44220
rect 15380 44040 15400 44200
rect 15580 44040 15600 44200
rect 15380 44020 15600 44040
rect 12644 39844 15100 39944
rect 12644 39108 12744 39844
rect 12644 38710 12656 39108
rect 12734 38710 12744 39108
rect 12644 38698 12744 38710
rect 12396 38638 13776 38658
rect 12396 38458 12536 38638
rect 12856 38458 12936 38638
rect 13356 38458 13776 38638
rect 12396 38438 13776 38458
rect 5156 38298 13776 38318
rect 5156 38118 5176 38298
rect 5476 38118 12716 38298
rect 12936 38118 13356 38298
rect 13576 38118 13776 38298
rect 5156 38098 13776 38118
rect 14536 38298 14656 38318
rect 14536 38078 14556 38298
rect 14636 38078 14656 38298
rect 14536 38058 14656 38078
rect 7426 37978 10676 37998
rect 7426 37818 7446 37978
rect 10656 37818 10676 37978
rect 14356 37838 14476 37858
rect 7426 37418 10676 37818
rect 12396 37818 14276 37838
rect 7426 37148 7436 37418
rect 10666 37148 10676 37418
rect 11576 37658 11836 37678
rect 11576 37178 11596 37658
rect 11816 37178 11836 37658
rect 12396 37638 12716 37818
rect 12936 37638 13356 37818
rect 13576 37638 13976 37818
rect 14256 37638 14276 37818
rect 12396 37618 14276 37638
rect 14356 37618 14376 37838
rect 14456 37618 14476 37838
rect 14356 37598 14476 37618
rect 11576 37158 11836 37178
rect 12396 37478 13776 37498
rect 12396 37298 12936 37478
rect 13356 37298 13496 37478
rect 12396 37178 13496 37298
rect 7426 37138 10676 37148
rect 7696 36988 7826 36998
rect 7696 36928 7706 36988
rect 7816 36928 7826 36988
rect 7696 36678 7826 36928
rect 7696 36608 7706 36678
rect 7816 36608 7826 36678
rect 7696 36598 7826 36608
rect 7856 36988 8186 36998
rect 7856 36768 7866 36988
rect 8136 36778 8186 36988
rect 7856 36618 8086 36768
rect 8176 36618 8186 36778
rect 7856 36598 8186 36618
rect 8216 36988 8346 36998
rect 8216 36918 8226 36988
rect 8336 36918 8346 36988
rect 8216 36668 8346 36918
rect 8216 36608 8226 36668
rect 8336 36608 8346 36668
rect 8216 36598 8346 36608
rect 8726 36988 8856 37008
rect 8726 36878 8736 36988
rect 8846 36878 8856 36988
rect 8726 36678 8856 36878
rect 8726 36608 8736 36678
rect 8846 36608 8856 36678
rect 8726 36598 8856 36608
rect 9246 36998 9376 37008
rect 9246 36918 9256 36998
rect 9366 36918 9376 36998
rect 9246 36668 9376 36918
rect 9246 36608 9256 36668
rect 9366 36608 9376 36668
rect 9246 36598 9376 36608
rect 9766 36998 9896 37008
rect 9766 36878 9776 36998
rect 9886 36878 9896 36998
rect 9766 36678 9896 36878
rect 10276 36998 10406 37008
rect 10276 36918 10286 36998
rect 10396 36918 10406 36998
rect 12396 36998 12936 37178
rect 13356 36998 13496 37178
rect 13676 36998 13776 37478
rect 12396 36978 13776 36998
rect 9766 36608 9776 36678
rect 9886 36608 9896 36678
rect 9946 36788 10246 36798
rect 9946 36618 9966 36788
rect 10236 36618 10246 36788
rect 9946 36608 10246 36618
rect 10276 36668 10406 36918
rect 10276 36608 10286 36668
rect 10396 36608 10406 36668
rect 11936 36838 13776 36858
rect 11936 36658 11956 36838
rect 12156 36658 12716 36838
rect 12936 36658 13356 36838
rect 13576 36658 13776 36838
rect 11936 36638 13776 36658
rect 14536 36838 14656 36858
rect 9766 36598 9896 36608
rect 10276 36598 10406 36608
rect 14536 36618 14556 36838
rect 14636 36618 14656 36838
rect 14536 36598 14656 36618
rect 7946 36558 10156 36568
rect 7946 36498 7966 36558
rect 8076 36498 8486 36558
rect 8596 36498 9006 36558
rect 9116 36498 9516 36558
rect 9626 36498 10026 36558
rect 10136 36498 10156 36558
rect 7946 36478 10156 36498
rect 6936 36368 9196 36408
rect 6936 36308 8946 36368
rect 9166 36308 9196 36368
rect 6936 36298 9196 36308
rect 6936 36128 7376 36298
rect 9266 36263 9626 36478
rect 14356 36378 14476 36398
rect 8476 36248 9626 36263
rect 8476 36173 8511 36248
rect 8566 36173 9541 36248
rect 9596 36173 9626 36248
rect 8476 36158 9626 36173
rect 12396 36358 14276 36378
rect 12396 36178 12716 36358
rect 12936 36178 13356 36358
rect 13576 36178 13976 36358
rect 14256 36178 14276 36358
rect 12396 36158 14276 36178
rect 14356 36158 14376 36378
rect 14456 36158 14476 36378
rect 14356 36138 14476 36158
rect 6936 36008 6946 36128
rect 7366 36008 7376 36128
rect 6936 35998 7376 36008
rect 7426 35848 7446 36098
rect 10656 35848 10676 36098
rect 7426 35678 10676 35848
rect 12396 36018 13776 36038
rect 12396 35838 12456 36018
rect 12856 35838 12936 36018
rect 13356 35838 13776 36018
rect 12396 35818 13776 35838
rect 7426 35518 7446 35678
rect 10656 35518 10676 35678
rect 7426 35498 10676 35518
rect 12456 35578 13576 35598
rect 12456 35478 12976 35578
rect 13356 35478 13576 35578
rect 12456 35418 12576 35478
rect 13536 35418 13576 35478
rect 12456 35398 13576 35418
rect 12196 35238 12416 35258
rect 12196 35058 12216 35238
rect 12396 35058 12416 35238
rect 12196 35038 12416 35058
rect 13476 35238 13696 35258
rect 13476 35058 13496 35238
rect 13676 35058 13696 35238
rect 13476 35038 13696 35058
rect 12456 34938 13576 34958
rect 12456 34778 12536 34938
rect 13556 34878 13576 34938
rect 12856 34778 13576 34878
rect 12456 34758 13576 34778
rect 15440 33936 15540 44020
rect 17080 44000 17320 44020
rect 17080 43820 17100 44000
rect 17300 43820 17320 44000
rect 17080 43800 17320 43820
rect 15760 43780 15980 43800
rect 15760 43620 15780 43780
rect 15960 43620 15980 43780
rect 15760 43600 15980 43620
rect 15820 38120 15920 43600
rect 16820 43540 17000 43560
rect 16820 43420 16840 43540
rect 16980 43420 17000 43540
rect 16820 43400 17000 43420
rect 16080 43340 16260 43360
rect 16080 43220 16100 43340
rect 16240 43220 16260 43340
rect 16080 43200 16260 43220
rect 12694 33836 15540 33936
rect 12694 33214 12794 33836
rect 12694 32886 12710 33214
rect 12782 32886 12794 33214
rect 12694 32870 12794 32886
rect 12416 32712 13796 32732
rect 12416 32532 12556 32712
rect 12876 32532 12956 32712
rect 13376 32532 13796 32712
rect 12416 32512 13796 32532
rect 5176 32372 13796 32392
rect 5176 32192 5196 32372
rect 5496 32192 12736 32372
rect 12956 32192 13376 32372
rect 13596 32192 13796 32372
rect 5176 32172 13796 32192
rect 14556 32372 14676 32392
rect 14556 32152 14576 32372
rect 14656 32152 14676 32372
rect 14556 32132 14676 32152
rect 7446 32052 10696 32072
rect 7446 31892 7466 32052
rect 10676 31892 10696 32052
rect 14376 31912 14496 31932
rect 7446 31492 10696 31892
rect 12416 31892 14296 31912
rect 7446 31222 7456 31492
rect 10686 31222 10696 31492
rect 11596 31732 11856 31752
rect 11596 31252 11616 31732
rect 11836 31252 11856 31732
rect 12416 31712 12736 31892
rect 12956 31712 13376 31892
rect 13596 31712 13996 31892
rect 14276 31712 14296 31892
rect 12416 31692 14296 31712
rect 14376 31692 14396 31912
rect 14476 31692 14496 31912
rect 14376 31672 14496 31692
rect 11596 31232 11856 31252
rect 12416 31552 13796 31572
rect 12416 31372 12956 31552
rect 13376 31372 13516 31552
rect 12416 31252 13516 31372
rect 7446 31212 10696 31222
rect 7716 31062 7846 31072
rect 7716 31002 7726 31062
rect 7836 31002 7846 31062
rect 7716 30752 7846 31002
rect 7716 30682 7726 30752
rect 7836 30682 7846 30752
rect 7716 30672 7846 30682
rect 7876 31062 8206 31072
rect 7876 30842 7886 31062
rect 8156 30852 8206 31062
rect 7876 30692 8106 30842
rect 8196 30692 8206 30852
rect 7876 30672 8206 30692
rect 8236 31062 8366 31072
rect 8236 30992 8246 31062
rect 8356 30992 8366 31062
rect 8236 30742 8366 30992
rect 8236 30682 8246 30742
rect 8356 30682 8366 30742
rect 8236 30672 8366 30682
rect 8746 31062 8876 31082
rect 8746 30952 8756 31062
rect 8866 30952 8876 31062
rect 8746 30752 8876 30952
rect 8746 30682 8756 30752
rect 8866 30682 8876 30752
rect 8746 30672 8876 30682
rect 9266 31072 9396 31082
rect 9266 30992 9276 31072
rect 9386 30992 9396 31072
rect 9266 30742 9396 30992
rect 9266 30682 9276 30742
rect 9386 30682 9396 30742
rect 9266 30672 9396 30682
rect 9786 31072 9916 31082
rect 9786 30952 9796 31072
rect 9906 30952 9916 31072
rect 9786 30752 9916 30952
rect 10296 31072 10426 31082
rect 10296 30992 10306 31072
rect 10416 30992 10426 31072
rect 12416 31072 12956 31252
rect 13376 31072 13516 31252
rect 13696 31072 13796 31552
rect 12416 31052 13796 31072
rect 9786 30682 9796 30752
rect 9906 30682 9916 30752
rect 9966 30862 10266 30872
rect 9966 30692 9986 30862
rect 10256 30692 10266 30862
rect 9966 30682 10266 30692
rect 10296 30742 10426 30992
rect 10296 30682 10306 30742
rect 10416 30682 10426 30742
rect 11956 30912 13796 30932
rect 11956 30732 11976 30912
rect 12176 30732 12736 30912
rect 12956 30732 13376 30912
rect 13596 30732 13796 30912
rect 11956 30712 13796 30732
rect 14556 30912 14676 30932
rect 9786 30672 9916 30682
rect 10296 30672 10426 30682
rect 14556 30692 14576 30912
rect 14656 30692 14676 30912
rect 14556 30672 14676 30692
rect 7966 30632 10176 30642
rect 7966 30572 7986 30632
rect 8096 30572 8506 30632
rect 8616 30572 9026 30632
rect 9136 30572 9536 30632
rect 9646 30572 10046 30632
rect 10156 30572 10176 30632
rect 7966 30552 10176 30572
rect 6956 30442 9216 30482
rect 6956 30382 8966 30442
rect 9186 30382 9216 30442
rect 6956 30372 9216 30382
rect 6956 30202 7396 30372
rect 9286 30337 9646 30552
rect 14376 30452 14496 30472
rect 8496 30322 9646 30337
rect 8496 30247 8531 30322
rect 8586 30247 9561 30322
rect 9616 30247 9646 30322
rect 8496 30232 9646 30247
rect 12416 30432 14296 30452
rect 12416 30252 12736 30432
rect 12956 30252 13376 30432
rect 13596 30252 13996 30432
rect 14276 30252 14296 30432
rect 12416 30232 14296 30252
rect 14376 30232 14396 30452
rect 14476 30232 14496 30452
rect 14376 30212 14496 30232
rect 6956 30082 6966 30202
rect 7386 30082 7396 30202
rect 6956 30072 7396 30082
rect 7446 29922 7466 30172
rect 10676 30132 11596 30172
rect 10676 29922 11456 30132
rect 7446 29752 11456 29922
rect 7446 29592 7466 29752
rect 10676 29692 11456 29752
rect 11556 29692 11596 30132
rect 12416 30092 13796 30112
rect 12416 29912 12476 30092
rect 12876 29912 12956 30092
rect 13376 29912 13796 30092
rect 12416 29892 13796 29912
rect 10676 29652 11596 29692
rect 12476 29652 13596 29672
rect 10676 29592 10696 29652
rect 7446 29572 10696 29592
rect 9536 29132 10696 29572
rect 12476 29552 12996 29652
rect 13376 29552 13596 29652
rect 12476 29492 12596 29552
rect 13556 29492 13596 29552
rect 12476 29472 13596 29492
rect 12216 29312 12436 29332
rect 9536 29052 9556 29132
rect 10676 29052 10696 29132
rect 9536 29012 10696 29052
rect 11616 29272 11816 29292
rect 11616 29012 11636 29272
rect 10836 28992 11636 29012
rect 10836 28812 10856 28992
rect 11796 28812 11816 29272
rect 12216 29132 12236 29312
rect 12416 29132 12436 29312
rect 12216 29112 12436 29132
rect 13496 29312 13716 29332
rect 13496 29132 13516 29312
rect 13696 29132 13716 29312
rect 13496 29112 13716 29132
rect 12476 29012 13596 29032
rect 12476 28852 12556 29012
rect 13576 28952 13596 29012
rect 12876 28852 13596 28952
rect 12476 28832 13596 28852
rect 10836 28792 11816 28812
rect 15821 27236 15920 38120
rect 12811 27137 15920 27236
rect 12811 26512 12910 27137
rect 12811 26080 12824 26512
rect 12898 26080 12910 26512
rect 12811 26067 12910 26080
rect 12536 26008 13916 26028
rect 12536 25828 12676 26008
rect 12996 25828 13076 26008
rect 13496 25828 13916 26008
rect 12536 25808 13916 25828
rect 5296 25668 13916 25688
rect 5296 25488 5316 25668
rect 5616 25488 12856 25668
rect 13076 25488 13496 25668
rect 13716 25488 13916 25668
rect 5296 25468 13916 25488
rect 14676 25668 14796 25688
rect 14676 25448 14696 25668
rect 14776 25448 14796 25668
rect 14676 25428 14796 25448
rect 7566 25348 10816 25368
rect 7566 25188 7586 25348
rect 10796 25188 10816 25348
rect 14496 25208 14616 25228
rect 7566 24788 10816 25188
rect 12536 25188 14416 25208
rect 7566 24518 7576 24788
rect 10806 24518 10816 24788
rect 11716 25028 11976 25048
rect 11716 24548 11736 25028
rect 11956 24548 11976 25028
rect 12536 25008 12856 25188
rect 13076 25008 13496 25188
rect 13716 25008 14116 25188
rect 14396 25008 14416 25188
rect 12536 24988 14416 25008
rect 14496 24988 14516 25208
rect 14596 24988 14616 25208
rect 14496 24968 14616 24988
rect 11716 24528 11976 24548
rect 12536 24848 13916 24868
rect 12536 24668 13076 24848
rect 13496 24668 13636 24848
rect 12536 24548 13636 24668
rect 7566 24508 10816 24518
rect 7836 24358 7966 24368
rect 7836 24298 7846 24358
rect 7956 24298 7966 24358
rect 7836 24048 7966 24298
rect 7836 23978 7846 24048
rect 7956 23978 7966 24048
rect 7836 23968 7966 23978
rect 7996 24358 8326 24368
rect 7996 24138 8006 24358
rect 8276 24148 8326 24358
rect 7996 23988 8226 24138
rect 8316 23988 8326 24148
rect 7996 23968 8326 23988
rect 8356 24358 8486 24368
rect 8356 24288 8366 24358
rect 8476 24288 8486 24358
rect 8356 24038 8486 24288
rect 8356 23978 8366 24038
rect 8476 23978 8486 24038
rect 8356 23968 8486 23978
rect 8866 24358 8996 24378
rect 8866 24248 8876 24358
rect 8986 24248 8996 24358
rect 8866 24048 8996 24248
rect 8866 23978 8876 24048
rect 8986 23978 8996 24048
rect 8866 23968 8996 23978
rect 9386 24368 9516 24378
rect 9386 24288 9396 24368
rect 9506 24288 9516 24368
rect 9386 24038 9516 24288
rect 9386 23978 9396 24038
rect 9506 23978 9516 24038
rect 9386 23968 9516 23978
rect 9906 24368 10036 24378
rect 9906 24248 9916 24368
rect 10026 24248 10036 24368
rect 9906 24048 10036 24248
rect 10416 24368 10546 24378
rect 10416 24288 10426 24368
rect 10536 24288 10546 24368
rect 12536 24368 13076 24548
rect 13496 24368 13636 24548
rect 13816 24368 13916 24848
rect 12536 24348 13916 24368
rect 9906 23978 9916 24048
rect 10026 23978 10036 24048
rect 10086 24158 10386 24168
rect 10086 23988 10106 24158
rect 10376 23988 10386 24158
rect 10086 23978 10386 23988
rect 10416 24038 10546 24288
rect 10416 23978 10426 24038
rect 10536 23978 10546 24038
rect 12076 24208 13916 24228
rect 12076 24028 12096 24208
rect 12296 24028 12856 24208
rect 13076 24028 13496 24208
rect 13716 24028 13916 24208
rect 12076 24008 13916 24028
rect 14676 24208 14796 24228
rect 9906 23968 10036 23978
rect 10416 23968 10546 23978
rect 14676 23988 14696 24208
rect 14776 23988 14796 24208
rect 14676 23968 14796 23988
rect 8086 23928 10296 23938
rect 8086 23868 8106 23928
rect 8216 23868 8626 23928
rect 8736 23868 9146 23928
rect 9256 23868 9656 23928
rect 9766 23868 10166 23928
rect 10276 23868 10296 23928
rect 8086 23848 10296 23868
rect 7076 23738 9336 23778
rect 7076 23678 9086 23738
rect 9306 23678 9336 23738
rect 7076 23668 9336 23678
rect 7076 23498 7516 23668
rect 9406 23633 9766 23848
rect 14496 23748 14616 23768
rect 8616 23618 9766 23633
rect 8616 23543 8651 23618
rect 8706 23543 9681 23618
rect 9736 23543 9766 23618
rect 8616 23528 9766 23543
rect 12536 23728 14416 23748
rect 12536 23548 12856 23728
rect 13076 23548 13496 23728
rect 13716 23548 14116 23728
rect 14396 23548 14416 23728
rect 12536 23528 14416 23548
rect 14496 23528 14516 23748
rect 14596 23528 14616 23748
rect 14496 23508 14616 23528
rect 7076 23378 7086 23498
rect 7506 23378 7516 23498
rect 7076 23368 7516 23378
rect 7566 23218 7586 23468
rect 10796 23428 11716 23468
rect 10796 23218 11576 23428
rect 7566 23048 11576 23218
rect 7566 22888 7586 23048
rect 10796 22988 11576 23048
rect 11676 22988 11716 23428
rect 12536 23388 13916 23408
rect 12536 23208 12596 23388
rect 12996 23208 13076 23388
rect 13496 23208 13916 23388
rect 12536 23188 13916 23208
rect 10796 22948 11716 22988
rect 12596 22948 13716 22968
rect 10796 22888 10816 22948
rect 7566 22868 10816 22888
rect 9656 22428 10816 22868
rect 12596 22848 13116 22948
rect 13496 22848 13716 22948
rect 12596 22788 12716 22848
rect 13676 22788 13716 22848
rect 12596 22768 13716 22788
rect 12336 22608 12556 22628
rect 9656 22348 9676 22428
rect 10796 22348 10816 22428
rect 9656 22308 10816 22348
rect 11736 22568 11936 22588
rect 11736 22308 11756 22568
rect 10956 22288 11756 22308
rect 10956 22108 10976 22288
rect 11916 22108 11936 22568
rect 12336 22428 12356 22608
rect 12536 22428 12556 22608
rect 12336 22408 12556 22428
rect 13616 22608 13836 22628
rect 13616 22428 13636 22608
rect 13816 22428 13836 22608
rect 13616 22408 13836 22428
rect 12596 22308 13716 22328
rect 12596 22148 12676 22308
rect 13696 22248 13716 22308
rect 12996 22148 13716 22248
rect 12596 22128 13716 22148
rect 10956 22088 11936 22108
rect 16120 20342 16220 43200
rect 16440 43140 16620 43160
rect 16440 43000 16460 43140
rect 16600 43000 16620 43140
rect 16440 42980 16620 43000
rect 12694 20242 16220 20342
rect 16480 20382 16580 42980
rect 16860 27300 16960 43400
rect 17140 34040 17240 43800
rect 17440 39824 17540 44260
rect 17440 39724 25516 39824
rect 25416 39258 25516 39724
rect 25416 38862 25432 39258
rect 25502 38862 25516 39258
rect 25416 38844 25516 38862
rect 25184 38756 26564 38776
rect 25184 38576 25324 38756
rect 25644 38576 25724 38756
rect 26144 38576 26564 38756
rect 25184 38556 26564 38576
rect 17944 38416 26564 38436
rect 17944 38236 17964 38416
rect 18264 38236 25504 38416
rect 25724 38236 26144 38416
rect 26364 38236 26564 38416
rect 17944 38216 26564 38236
rect 27324 38416 27444 38436
rect 27324 38196 27344 38416
rect 27424 38196 27444 38416
rect 27324 38176 27444 38196
rect 20214 38096 23464 38116
rect 20214 37936 20234 38096
rect 23444 37936 23464 38096
rect 27144 37956 27264 37976
rect 20214 37536 23464 37936
rect 25184 37936 27064 37956
rect 20214 37266 20224 37536
rect 23454 37266 23464 37536
rect 24364 37776 24624 37796
rect 24364 37296 24384 37776
rect 24604 37296 24624 37776
rect 25184 37756 25504 37936
rect 25724 37756 26144 37936
rect 26364 37756 26764 37936
rect 27044 37756 27064 37936
rect 25184 37736 27064 37756
rect 27144 37736 27164 37956
rect 27244 37736 27264 37956
rect 27144 37716 27264 37736
rect 24364 37276 24624 37296
rect 25184 37596 26564 37616
rect 25184 37416 25724 37596
rect 26144 37416 26284 37596
rect 25184 37296 26284 37416
rect 20214 37256 23464 37266
rect 20484 37106 20614 37116
rect 20484 37046 20494 37106
rect 20604 37046 20614 37106
rect 20484 36796 20614 37046
rect 20484 36726 20494 36796
rect 20604 36726 20614 36796
rect 20484 36716 20614 36726
rect 20644 37106 20974 37116
rect 20644 36886 20654 37106
rect 20924 36896 20974 37106
rect 20644 36736 20874 36886
rect 20964 36736 20974 36896
rect 20644 36716 20974 36736
rect 21004 37106 21134 37116
rect 21004 37036 21014 37106
rect 21124 37036 21134 37106
rect 21004 36786 21134 37036
rect 21004 36726 21014 36786
rect 21124 36726 21134 36786
rect 21004 36716 21134 36726
rect 21514 37106 21644 37126
rect 21514 36996 21524 37106
rect 21634 36996 21644 37106
rect 21514 36796 21644 36996
rect 21514 36726 21524 36796
rect 21634 36726 21644 36796
rect 21514 36716 21644 36726
rect 22034 37116 22164 37126
rect 22034 37036 22044 37116
rect 22154 37036 22164 37116
rect 22034 36786 22164 37036
rect 22034 36726 22044 36786
rect 22154 36726 22164 36786
rect 22034 36716 22164 36726
rect 22554 37116 22684 37126
rect 22554 36996 22564 37116
rect 22674 36996 22684 37116
rect 22554 36796 22684 36996
rect 23064 37116 23194 37126
rect 23064 37036 23074 37116
rect 23184 37036 23194 37116
rect 25184 37116 25724 37296
rect 26144 37116 26284 37296
rect 26464 37116 26564 37596
rect 25184 37096 26564 37116
rect 22554 36726 22564 36796
rect 22674 36726 22684 36796
rect 22734 36906 23034 36916
rect 22734 36736 22754 36906
rect 23024 36736 23034 36906
rect 22734 36726 23034 36736
rect 23064 36786 23194 37036
rect 23064 36726 23074 36786
rect 23184 36726 23194 36786
rect 24724 36956 26564 36976
rect 24724 36776 24744 36956
rect 24944 36776 25504 36956
rect 25724 36776 26144 36956
rect 26364 36776 26564 36956
rect 24724 36756 26564 36776
rect 27324 36956 27444 36976
rect 22554 36716 22684 36726
rect 23064 36716 23194 36726
rect 27324 36736 27344 36956
rect 27424 36736 27444 36956
rect 27324 36716 27444 36736
rect 20734 36676 22944 36686
rect 20734 36616 20754 36676
rect 20864 36616 21274 36676
rect 21384 36616 21794 36676
rect 21904 36616 22304 36676
rect 22414 36616 22814 36676
rect 22924 36616 22944 36676
rect 20734 36596 22944 36616
rect 19724 36486 21984 36526
rect 19724 36426 21734 36486
rect 21954 36426 21984 36486
rect 19724 36416 21984 36426
rect 19724 36246 20164 36416
rect 22054 36381 22414 36596
rect 27144 36496 27264 36516
rect 21264 36366 22414 36381
rect 21264 36291 21299 36366
rect 21354 36291 22329 36366
rect 22384 36291 22414 36366
rect 21264 36276 22414 36291
rect 25184 36476 27064 36496
rect 25184 36296 25504 36476
rect 25724 36296 26144 36476
rect 26364 36296 26764 36476
rect 27044 36296 27064 36476
rect 25184 36276 27064 36296
rect 27144 36276 27164 36496
rect 27244 36276 27264 36496
rect 27144 36256 27264 36276
rect 19724 36126 19734 36246
rect 20154 36126 20164 36246
rect 19724 36116 20164 36126
rect 20214 35966 20234 36216
rect 23444 36176 24364 36216
rect 23444 35966 24224 36176
rect 20214 35796 24224 35966
rect 20214 35636 20234 35796
rect 23444 35736 24224 35796
rect 24324 35736 24364 36176
rect 25184 36136 26564 36156
rect 25184 35956 25244 36136
rect 25644 35956 25724 36136
rect 26144 35956 26564 36136
rect 25184 35936 26564 35956
rect 23444 35696 24364 35736
rect 25244 35696 26364 35716
rect 23444 35636 23464 35696
rect 20214 35616 23464 35636
rect 22304 35176 23464 35616
rect 25244 35596 25764 35696
rect 26144 35596 26364 35696
rect 25244 35536 25364 35596
rect 26324 35536 26364 35596
rect 25244 35516 26364 35536
rect 24984 35356 25204 35376
rect 22304 35096 22324 35176
rect 23444 35096 23464 35176
rect 22304 35056 23464 35096
rect 24384 35316 24584 35336
rect 24384 35056 24404 35316
rect 23604 35036 24404 35056
rect 23604 34856 23624 35036
rect 24564 34856 24584 35316
rect 24984 35176 25004 35356
rect 25184 35176 25204 35356
rect 24984 35156 25204 35176
rect 26264 35356 26484 35376
rect 26264 35176 26284 35356
rect 26464 35176 26484 35356
rect 26264 35156 26484 35176
rect 25244 35056 26364 35076
rect 25244 34896 25324 35056
rect 26344 34996 26364 35056
rect 25644 34896 26364 34996
rect 25244 34876 26364 34896
rect 23604 34836 24584 34856
rect 17140 33940 25422 34040
rect 25322 33132 25422 33940
rect 25322 32804 25336 33132
rect 25408 32804 25422 33132
rect 25322 32792 25422 32804
rect 25148 32636 26528 32656
rect 25148 32456 25288 32636
rect 25608 32456 25688 32636
rect 26108 32456 26528 32636
rect 25148 32436 26528 32456
rect 17908 32296 26528 32316
rect 17908 32116 17928 32296
rect 18228 32116 25468 32296
rect 25688 32116 26108 32296
rect 26328 32116 26528 32296
rect 17908 32096 26528 32116
rect 27288 32296 27408 32316
rect 27288 32076 27308 32296
rect 27388 32076 27408 32296
rect 27288 32056 27408 32076
rect 20178 31976 23428 31996
rect 20178 31816 20198 31976
rect 23408 31816 23428 31976
rect 27108 31836 27228 31856
rect 20178 31416 23428 31816
rect 25148 31816 27028 31836
rect 20178 31146 20188 31416
rect 23418 31146 23428 31416
rect 24328 31656 24588 31676
rect 24328 31176 24348 31656
rect 24568 31176 24588 31656
rect 25148 31636 25468 31816
rect 25688 31636 26108 31816
rect 26328 31636 26728 31816
rect 27008 31636 27028 31816
rect 25148 31616 27028 31636
rect 27108 31616 27128 31836
rect 27208 31616 27228 31836
rect 27108 31596 27228 31616
rect 24328 31156 24588 31176
rect 25148 31476 26528 31496
rect 25148 31296 25688 31476
rect 26108 31296 26248 31476
rect 25148 31176 26248 31296
rect 20178 31136 23428 31146
rect 20448 30986 20578 30996
rect 20448 30926 20458 30986
rect 20568 30926 20578 30986
rect 20448 30676 20578 30926
rect 20448 30606 20458 30676
rect 20568 30606 20578 30676
rect 20448 30596 20578 30606
rect 20608 30986 20938 30996
rect 20608 30766 20618 30986
rect 20888 30776 20938 30986
rect 20608 30616 20838 30766
rect 20928 30616 20938 30776
rect 20608 30596 20938 30616
rect 20968 30986 21098 30996
rect 20968 30916 20978 30986
rect 21088 30916 21098 30986
rect 20968 30666 21098 30916
rect 20968 30606 20978 30666
rect 21088 30606 21098 30666
rect 20968 30596 21098 30606
rect 21478 30986 21608 31006
rect 21478 30876 21488 30986
rect 21598 30876 21608 30986
rect 21478 30676 21608 30876
rect 21478 30606 21488 30676
rect 21598 30606 21608 30676
rect 21478 30596 21608 30606
rect 21998 30996 22128 31006
rect 21998 30916 22008 30996
rect 22118 30916 22128 30996
rect 21998 30666 22128 30916
rect 21998 30606 22008 30666
rect 22118 30606 22128 30666
rect 21998 30596 22128 30606
rect 22518 30996 22648 31006
rect 22518 30876 22528 30996
rect 22638 30876 22648 30996
rect 22518 30676 22648 30876
rect 23028 30996 23158 31006
rect 23028 30916 23038 30996
rect 23148 30916 23158 30996
rect 25148 30996 25688 31176
rect 26108 30996 26248 31176
rect 26428 30996 26528 31476
rect 25148 30976 26528 30996
rect 22518 30606 22528 30676
rect 22638 30606 22648 30676
rect 22698 30786 22998 30796
rect 22698 30616 22718 30786
rect 22988 30616 22998 30786
rect 22698 30606 22998 30616
rect 23028 30666 23158 30916
rect 23028 30606 23038 30666
rect 23148 30606 23158 30666
rect 24688 30836 26528 30856
rect 24688 30656 24708 30836
rect 24908 30656 25468 30836
rect 25688 30656 26108 30836
rect 26328 30656 26528 30836
rect 24688 30636 26528 30656
rect 27288 30836 27408 30856
rect 22518 30596 22648 30606
rect 23028 30596 23158 30606
rect 27288 30616 27308 30836
rect 27388 30616 27408 30836
rect 27288 30596 27408 30616
rect 20698 30556 22908 30566
rect 20698 30496 20718 30556
rect 20828 30496 21238 30556
rect 21348 30496 21758 30556
rect 21868 30496 22268 30556
rect 22378 30496 22778 30556
rect 22888 30496 22908 30556
rect 20698 30476 22908 30496
rect 19688 30366 21948 30406
rect 19688 30306 21698 30366
rect 21918 30306 21948 30366
rect 19688 30296 21948 30306
rect 19688 30126 20128 30296
rect 22018 30261 22378 30476
rect 27108 30376 27228 30396
rect 21228 30246 22378 30261
rect 21228 30171 21263 30246
rect 21318 30171 22293 30246
rect 22348 30171 22378 30246
rect 21228 30156 22378 30171
rect 25148 30356 27028 30376
rect 25148 30176 25468 30356
rect 25688 30176 26108 30356
rect 26328 30176 26728 30356
rect 27008 30176 27028 30356
rect 25148 30156 27028 30176
rect 27108 30156 27128 30376
rect 27208 30156 27228 30376
rect 27108 30136 27228 30156
rect 19688 30006 19698 30126
rect 20118 30006 20128 30126
rect 19688 29996 20128 30006
rect 20178 29846 20198 30096
rect 23408 30056 24328 30096
rect 23408 29846 24188 30056
rect 20178 29676 24188 29846
rect 20178 29516 20198 29676
rect 23408 29616 24188 29676
rect 24288 29616 24328 30056
rect 25148 30016 26528 30036
rect 25148 29836 25208 30016
rect 25608 29836 25688 30016
rect 26108 29836 26528 30016
rect 25148 29816 26528 29836
rect 23408 29576 24328 29616
rect 25208 29576 26328 29596
rect 23408 29516 23428 29576
rect 20178 29496 23428 29516
rect 22268 29056 23428 29496
rect 25208 29476 25728 29576
rect 26108 29476 26328 29576
rect 25208 29416 25328 29476
rect 26288 29416 26328 29476
rect 25208 29396 26328 29416
rect 24948 29236 25168 29256
rect 22268 28976 22288 29056
rect 23408 28976 23428 29056
rect 22268 28936 23428 28976
rect 24348 29196 24548 29216
rect 24348 28936 24368 29196
rect 23568 28916 24368 28936
rect 23568 28736 23588 28916
rect 24528 28736 24548 29196
rect 24948 29056 24968 29236
rect 25148 29056 25168 29236
rect 24948 29036 25168 29056
rect 26228 29236 26448 29256
rect 26228 29056 26248 29236
rect 26428 29056 26448 29236
rect 26228 29036 26448 29056
rect 25208 28936 26328 28956
rect 25208 28776 25288 28936
rect 26308 28876 26328 28936
rect 25608 28776 26328 28876
rect 25208 28756 26328 28776
rect 23568 28716 24548 28736
rect 16860 27200 25602 27300
rect 16860 27174 16960 27200
rect 25502 26382 25602 27200
rect 25502 25988 25518 26382
rect 25586 25988 25602 26382
rect 25502 25970 25602 25988
rect 25244 25878 26624 25898
rect 25244 25698 25384 25878
rect 25704 25698 25784 25878
rect 26204 25698 26624 25878
rect 25244 25678 26624 25698
rect 18004 25538 26624 25558
rect 18004 25358 18024 25538
rect 18324 25358 25564 25538
rect 25784 25358 26204 25538
rect 26424 25358 26624 25538
rect 18004 25338 26624 25358
rect 27384 25538 27504 25558
rect 27384 25318 27404 25538
rect 27484 25318 27504 25538
rect 27384 25298 27504 25318
rect 20274 25218 23524 25238
rect 20274 25058 20294 25218
rect 23504 25058 23524 25218
rect 27204 25078 27324 25098
rect 20274 24658 23524 25058
rect 25244 25058 27124 25078
rect 20274 24388 20284 24658
rect 23514 24388 23524 24658
rect 24424 24898 24684 24918
rect 24424 24418 24444 24898
rect 24664 24418 24684 24898
rect 25244 24878 25564 25058
rect 25784 24878 26204 25058
rect 26424 24878 26824 25058
rect 27104 24878 27124 25058
rect 25244 24858 27124 24878
rect 27204 24858 27224 25078
rect 27304 24858 27324 25078
rect 27204 24838 27324 24858
rect 24424 24398 24684 24418
rect 25244 24718 26624 24738
rect 25244 24538 25784 24718
rect 26204 24538 26344 24718
rect 25244 24418 26344 24538
rect 20274 24378 23524 24388
rect 20544 24228 20674 24238
rect 20544 24168 20554 24228
rect 20664 24168 20674 24228
rect 20544 23918 20674 24168
rect 20544 23848 20554 23918
rect 20664 23848 20674 23918
rect 20544 23838 20674 23848
rect 20704 24228 21034 24238
rect 20704 24008 20714 24228
rect 20984 24018 21034 24228
rect 20704 23858 20934 24008
rect 21024 23858 21034 24018
rect 20704 23838 21034 23858
rect 21064 24228 21194 24238
rect 21064 24158 21074 24228
rect 21184 24158 21194 24228
rect 21064 23908 21194 24158
rect 21064 23848 21074 23908
rect 21184 23848 21194 23908
rect 21064 23838 21194 23848
rect 21574 24228 21704 24248
rect 21574 24118 21584 24228
rect 21694 24118 21704 24228
rect 21574 23918 21704 24118
rect 21574 23848 21584 23918
rect 21694 23848 21704 23918
rect 21574 23838 21704 23848
rect 22094 24238 22224 24248
rect 22094 24158 22104 24238
rect 22214 24158 22224 24238
rect 22094 23908 22224 24158
rect 22094 23848 22104 23908
rect 22214 23848 22224 23908
rect 22094 23838 22224 23848
rect 22614 24238 22744 24248
rect 22614 24118 22624 24238
rect 22734 24118 22744 24238
rect 22614 23918 22744 24118
rect 23124 24238 23254 24248
rect 23124 24158 23134 24238
rect 23244 24158 23254 24238
rect 25244 24238 25784 24418
rect 26204 24238 26344 24418
rect 26524 24238 26624 24718
rect 25244 24218 26624 24238
rect 22614 23848 22624 23918
rect 22734 23848 22744 23918
rect 22794 24028 23094 24038
rect 22794 23858 22814 24028
rect 23084 23858 23094 24028
rect 22794 23848 23094 23858
rect 23124 23908 23254 24158
rect 23124 23848 23134 23908
rect 23244 23848 23254 23908
rect 24784 24078 26624 24098
rect 24784 23898 24804 24078
rect 25004 23898 25564 24078
rect 25784 23898 26204 24078
rect 26424 23898 26624 24078
rect 24784 23878 26624 23898
rect 27384 24078 27504 24098
rect 22614 23838 22744 23848
rect 23124 23838 23254 23848
rect 27384 23858 27404 24078
rect 27484 23858 27504 24078
rect 27384 23838 27504 23858
rect 20794 23798 23004 23808
rect 20794 23738 20814 23798
rect 20924 23738 21334 23798
rect 21444 23738 21854 23798
rect 21964 23738 22364 23798
rect 22474 23738 22874 23798
rect 22984 23738 23004 23798
rect 20794 23718 23004 23738
rect 19784 23608 22044 23648
rect 19784 23548 21794 23608
rect 22014 23548 22044 23608
rect 19784 23538 22044 23548
rect 19784 23368 20224 23538
rect 22114 23503 22474 23718
rect 27204 23618 27324 23638
rect 21324 23488 22474 23503
rect 21324 23413 21359 23488
rect 21414 23413 22389 23488
rect 22444 23413 22474 23488
rect 21324 23398 22474 23413
rect 25244 23598 27124 23618
rect 25244 23418 25564 23598
rect 25784 23418 26204 23598
rect 26424 23418 26824 23598
rect 27104 23418 27124 23598
rect 25244 23398 27124 23418
rect 27204 23398 27224 23618
rect 27304 23398 27324 23618
rect 27204 23378 27324 23398
rect 19784 23248 19794 23368
rect 20214 23248 20224 23368
rect 19784 23238 20224 23248
rect 20274 23088 20294 23338
rect 23504 23298 24424 23338
rect 23504 23088 24284 23298
rect 20274 22918 24284 23088
rect 20274 22758 20294 22918
rect 23504 22858 24284 22918
rect 24384 22858 24424 23298
rect 25244 23258 26624 23278
rect 25244 23078 25304 23258
rect 25704 23078 25784 23258
rect 26204 23078 26624 23258
rect 25244 23058 26624 23078
rect 23504 22818 24424 22858
rect 25304 22818 26424 22838
rect 23504 22758 23524 22818
rect 20274 22738 23524 22758
rect 22364 22298 23524 22738
rect 25304 22718 25824 22818
rect 26204 22718 26424 22818
rect 25304 22658 25424 22718
rect 26384 22658 26424 22718
rect 25304 22638 26424 22658
rect 25044 22478 25264 22498
rect 22364 22218 22384 22298
rect 23504 22218 23524 22298
rect 22364 22178 23524 22218
rect 24444 22438 24644 22458
rect 24444 22178 24464 22438
rect 23664 22158 24464 22178
rect 23664 21978 23684 22158
rect 24624 21978 24644 22438
rect 25044 22298 25064 22478
rect 25244 22298 25264 22478
rect 25044 22278 25264 22298
rect 26324 22478 26544 22498
rect 26324 22298 26344 22478
rect 26524 22298 26544 22478
rect 26324 22278 26544 22298
rect 25304 22178 26424 22198
rect 25304 22018 25384 22178
rect 26404 22118 26424 22178
rect 25704 22018 26424 22118
rect 25304 21998 26424 22018
rect 23664 21958 24644 21978
rect 16480 20282 25938 20382
rect 12694 19464 12794 20242
rect 12694 19126 12706 19464
rect 12780 19126 12794 19464
rect 12694 19108 12794 19126
rect 25838 19334 25938 20282
rect 12412 18962 13792 18982
rect 12412 18782 12552 18962
rect 12872 18782 12952 18962
rect 13372 18782 13792 18962
rect 25838 18942 25852 19334
rect 25926 18942 25938 19334
rect 25838 18928 25938 18942
rect 12412 18762 13792 18782
rect 25594 18832 26974 18852
rect 25594 18652 25734 18832
rect 26054 18652 26134 18832
rect 26554 18652 26974 18832
rect 5172 18622 13792 18642
rect 5172 18442 5192 18622
rect 5492 18442 12732 18622
rect 12952 18442 13372 18622
rect 13592 18442 13792 18622
rect 5172 18422 13792 18442
rect 14552 18622 14672 18642
rect 25594 18632 26974 18652
rect 14552 18402 14572 18622
rect 14652 18402 14672 18622
rect 14552 18382 14672 18402
rect 18354 18492 26974 18512
rect 7442 18302 10692 18322
rect 7442 18142 7462 18302
rect 10672 18142 10692 18302
rect 18354 18312 18374 18492
rect 18674 18312 25914 18492
rect 26134 18312 26554 18492
rect 26774 18312 26974 18492
rect 18354 18292 26974 18312
rect 27734 18492 27854 18512
rect 27734 18272 27754 18492
rect 27834 18272 27854 18492
rect 27734 18252 27854 18272
rect 14372 18162 14492 18182
rect 7442 17742 10692 18142
rect 12412 18142 14292 18162
rect 7442 17472 7452 17742
rect 10682 17472 10692 17742
rect 11592 17982 11852 18002
rect 11592 17502 11612 17982
rect 11832 17502 11852 17982
rect 12412 17962 12732 18142
rect 12952 17962 13372 18142
rect 13592 17962 13992 18142
rect 14272 17962 14292 18142
rect 12412 17942 14292 17962
rect 14372 17942 14392 18162
rect 14472 17942 14492 18162
rect 14372 17922 14492 17942
rect 20624 18172 23874 18192
rect 20624 18012 20644 18172
rect 23854 18012 23874 18172
rect 27554 18032 27674 18052
rect 11592 17482 11852 17502
rect 12412 17802 13792 17822
rect 12412 17622 12952 17802
rect 13372 17622 13512 17802
rect 12412 17502 13512 17622
rect 7442 17462 10692 17472
rect 7712 17312 7842 17322
rect 7712 17252 7722 17312
rect 7832 17252 7842 17312
rect 7712 17002 7842 17252
rect 7712 16932 7722 17002
rect 7832 16932 7842 17002
rect 7712 16922 7842 16932
rect 7872 17312 8202 17322
rect 7872 17092 7882 17312
rect 8152 17102 8202 17312
rect 7872 16942 8102 17092
rect 8192 16942 8202 17102
rect 7872 16922 8202 16942
rect 8232 17312 8362 17322
rect 8232 17242 8242 17312
rect 8352 17242 8362 17312
rect 8232 16992 8362 17242
rect 8232 16932 8242 16992
rect 8352 16932 8362 16992
rect 8232 16922 8362 16932
rect 8742 17312 8872 17332
rect 8742 17202 8752 17312
rect 8862 17202 8872 17312
rect 8742 17002 8872 17202
rect 8742 16932 8752 17002
rect 8862 16932 8872 17002
rect 8742 16922 8872 16932
rect 9262 17322 9392 17332
rect 9262 17242 9272 17322
rect 9382 17242 9392 17322
rect 9262 16992 9392 17242
rect 9262 16932 9272 16992
rect 9382 16932 9392 16992
rect 9262 16922 9392 16932
rect 9782 17322 9912 17332
rect 9782 17202 9792 17322
rect 9902 17202 9912 17322
rect 9782 17002 9912 17202
rect 10292 17322 10422 17332
rect 10292 17242 10302 17322
rect 10412 17242 10422 17322
rect 12412 17322 12952 17502
rect 13372 17322 13512 17502
rect 13692 17322 13792 17802
rect 20624 17612 23874 18012
rect 25594 18012 27474 18032
rect 20624 17342 20634 17612
rect 23864 17342 23874 17612
rect 24774 17852 25034 17872
rect 24774 17372 24794 17852
rect 25014 17372 25034 17852
rect 25594 17832 25914 18012
rect 26134 17832 26554 18012
rect 26774 17832 27174 18012
rect 27454 17832 27474 18012
rect 25594 17812 27474 17832
rect 27554 17812 27574 18032
rect 27654 17812 27674 18032
rect 27554 17792 27674 17812
rect 24774 17352 25034 17372
rect 25594 17672 26974 17692
rect 25594 17492 26134 17672
rect 26554 17492 26694 17672
rect 25594 17372 26694 17492
rect 20624 17332 23874 17342
rect 12412 17302 13792 17322
rect 9782 16932 9792 17002
rect 9902 16932 9912 17002
rect 9962 17112 10262 17122
rect 9962 16942 9982 17112
rect 10252 16942 10262 17112
rect 9962 16932 10262 16942
rect 10292 16992 10422 17242
rect 20894 17182 21024 17192
rect 10292 16932 10302 16992
rect 10412 16932 10422 16992
rect 11952 17162 13792 17182
rect 11952 16982 11972 17162
rect 12172 16982 12732 17162
rect 12952 16982 13372 17162
rect 13592 16982 13792 17162
rect 11952 16962 13792 16982
rect 14552 17162 14672 17182
rect 9782 16922 9912 16932
rect 10292 16922 10422 16932
rect 14552 16942 14572 17162
rect 14652 16942 14672 17162
rect 14552 16922 14672 16942
rect 20894 17122 20904 17182
rect 21014 17122 21024 17182
rect 7962 16882 10172 16892
rect 7962 16822 7982 16882
rect 8092 16822 8502 16882
rect 8612 16822 9022 16882
rect 9132 16822 9532 16882
rect 9642 16822 10042 16882
rect 10152 16822 10172 16882
rect 7962 16802 10172 16822
rect 20894 16872 21024 17122
rect 20894 16802 20904 16872
rect 21014 16802 21024 16872
rect 6952 16692 9212 16732
rect 6952 16632 8962 16692
rect 9182 16632 9212 16692
rect 6952 16622 9212 16632
rect 6952 16452 7392 16622
rect 9282 16587 9642 16802
rect 20894 16792 21024 16802
rect 21054 17182 21384 17192
rect 21054 16962 21064 17182
rect 21334 16972 21384 17182
rect 21054 16812 21284 16962
rect 21374 16812 21384 16972
rect 21054 16792 21384 16812
rect 21414 17182 21544 17192
rect 21414 17112 21424 17182
rect 21534 17112 21544 17182
rect 21414 16862 21544 17112
rect 21414 16802 21424 16862
rect 21534 16802 21544 16862
rect 21414 16792 21544 16802
rect 21924 17182 22054 17202
rect 21924 17072 21934 17182
rect 22044 17072 22054 17182
rect 21924 16872 22054 17072
rect 21924 16802 21934 16872
rect 22044 16802 22054 16872
rect 21924 16792 22054 16802
rect 22444 17192 22574 17202
rect 22444 17112 22454 17192
rect 22564 17112 22574 17192
rect 22444 16862 22574 17112
rect 22444 16802 22454 16862
rect 22564 16802 22574 16862
rect 22444 16792 22574 16802
rect 22964 17192 23094 17202
rect 22964 17072 22974 17192
rect 23084 17072 23094 17192
rect 22964 16872 23094 17072
rect 23474 17192 23604 17202
rect 23474 17112 23484 17192
rect 23594 17112 23604 17192
rect 25594 17192 26134 17372
rect 26554 17192 26694 17372
rect 26874 17192 26974 17672
rect 25594 17172 26974 17192
rect 22964 16802 22974 16872
rect 23084 16802 23094 16872
rect 23144 16982 23444 16992
rect 23144 16812 23164 16982
rect 23434 16812 23444 16982
rect 23144 16802 23444 16812
rect 23474 16862 23604 17112
rect 23474 16802 23484 16862
rect 23594 16802 23604 16862
rect 25134 17032 26974 17052
rect 25134 16852 25154 17032
rect 25354 16852 25914 17032
rect 26134 16852 26554 17032
rect 26774 16852 26974 17032
rect 25134 16832 26974 16852
rect 27734 17032 27854 17052
rect 22964 16792 23094 16802
rect 23474 16792 23604 16802
rect 27734 16812 27754 17032
rect 27834 16812 27854 17032
rect 27734 16792 27854 16812
rect 21144 16752 23354 16762
rect 14372 16702 14492 16722
rect 8492 16572 9642 16587
rect 8492 16497 8527 16572
rect 8582 16497 9557 16572
rect 9612 16497 9642 16572
rect 8492 16482 9642 16497
rect 12412 16682 14292 16702
rect 12412 16502 12732 16682
rect 12952 16502 13372 16682
rect 13592 16502 13992 16682
rect 14272 16502 14292 16682
rect 12412 16482 14292 16502
rect 14372 16482 14392 16702
rect 14472 16482 14492 16702
rect 21144 16692 21164 16752
rect 21274 16692 21684 16752
rect 21794 16692 22204 16752
rect 22314 16692 22714 16752
rect 22824 16692 23224 16752
rect 23334 16692 23354 16752
rect 21144 16672 23354 16692
rect 14372 16462 14492 16482
rect 20134 16562 22394 16602
rect 20134 16502 22144 16562
rect 22364 16502 22394 16562
rect 20134 16492 22394 16502
rect 6952 16332 6962 16452
rect 7382 16332 7392 16452
rect 6952 16322 7392 16332
rect 7442 16172 7462 16422
rect 10672 16382 11592 16422
rect 10672 16172 11452 16382
rect 7442 16002 11452 16172
rect 7442 15842 7462 16002
rect 10672 15942 11452 16002
rect 11552 15942 11592 16382
rect 12412 16342 13792 16362
rect 12412 16162 12472 16342
rect 12872 16162 12952 16342
rect 13372 16162 13792 16342
rect 20134 16322 20574 16492
rect 22464 16457 22824 16672
rect 27554 16572 27674 16592
rect 21674 16442 22824 16457
rect 21674 16367 21709 16442
rect 21764 16367 22739 16442
rect 22794 16367 22824 16442
rect 21674 16352 22824 16367
rect 25594 16552 27474 16572
rect 25594 16372 25914 16552
rect 26134 16372 26554 16552
rect 26774 16372 27174 16552
rect 27454 16372 27474 16552
rect 25594 16352 27474 16372
rect 27554 16352 27574 16572
rect 27654 16352 27674 16572
rect 27554 16332 27674 16352
rect 20134 16202 20144 16322
rect 20564 16202 20574 16322
rect 20134 16192 20574 16202
rect 12412 16142 13792 16162
rect 10672 15902 11592 15942
rect 20624 16042 20644 16292
rect 23854 16252 24774 16292
rect 23854 16042 24634 16252
rect 12472 15902 13592 15922
rect 10672 15842 10692 15902
rect 7442 15822 10692 15842
rect 9532 15382 10692 15822
rect 12472 15802 12992 15902
rect 13372 15802 13592 15902
rect 12472 15742 12592 15802
rect 13552 15742 13592 15802
rect 12472 15722 13592 15742
rect 20624 15872 24634 16042
rect 20624 15712 20644 15872
rect 23854 15812 24634 15872
rect 24734 15812 24774 16252
rect 25594 16212 26974 16232
rect 25594 16032 25654 16212
rect 26054 16032 26134 16212
rect 26554 16032 26974 16212
rect 25594 16012 26974 16032
rect 23854 15772 24774 15812
rect 25654 15772 26774 15792
rect 23854 15712 23874 15772
rect 20624 15692 23874 15712
rect 12212 15562 12432 15582
rect 9532 15302 9552 15382
rect 10672 15302 10692 15382
rect 9532 15262 10692 15302
rect 11612 15522 11812 15542
rect 11612 15262 11632 15522
rect 10832 15242 11632 15262
rect 10832 15062 10852 15242
rect 11792 15062 11812 15522
rect 12212 15382 12232 15562
rect 12412 15382 12432 15562
rect 12212 15362 12432 15382
rect 13492 15562 13712 15582
rect 13492 15382 13512 15562
rect 13692 15382 13712 15562
rect 13492 15362 13712 15382
rect 12472 15262 13592 15282
rect 12472 15102 12552 15262
rect 13572 15202 13592 15262
rect 12872 15102 13592 15202
rect 22714 15252 23874 15692
rect 25654 15672 26174 15772
rect 26554 15672 26774 15772
rect 25654 15612 25774 15672
rect 26734 15612 26774 15672
rect 25654 15592 26774 15612
rect 25394 15432 25614 15452
rect 22714 15172 22734 15252
rect 23854 15172 23874 15252
rect 22714 15132 23874 15172
rect 24794 15392 24994 15412
rect 24794 15132 24814 15392
rect 12472 15082 13592 15102
rect 24014 15112 24814 15132
rect 10832 15042 11812 15062
rect 24014 14932 24034 15112
rect 24974 14932 24994 15392
rect 25394 15252 25414 15432
rect 25594 15252 25614 15432
rect 25394 15232 25614 15252
rect 26674 15432 26894 15452
rect 26674 15252 26694 15432
rect 26874 15252 26894 15432
rect 26674 15232 26894 15252
rect 25654 15132 26774 15152
rect 25654 14972 25734 15132
rect 26754 15072 26774 15132
rect 26054 14972 26774 15072
rect 25654 14952 26774 14972
rect 24014 14912 24994 14932
<< via2 >>
rect 14980 44480 15120 44600
rect 17400 44280 17580 44400
rect 15400 44040 15580 44200
rect 12656 38710 12734 39108
rect 12536 38458 12856 38638
rect 5176 38118 5476 38298
rect 14556 38078 14636 38298
rect 7436 37258 10666 37418
rect 7436 37178 7446 37258
rect 7446 37178 10606 37258
rect 10606 37178 10666 37258
rect 7436 37148 10666 37178
rect 11596 37178 11816 37658
rect 13976 37638 14256 37818
rect 14376 37618 14456 37838
rect 7706 36668 7816 36678
rect 7706 36608 7816 36668
rect 7866 36778 8136 36988
rect 7866 36768 8086 36778
rect 8086 36768 8136 36778
rect 8226 36928 8336 36988
rect 8226 36918 8336 36928
rect 8736 36668 8846 36678
rect 8736 36608 8846 36668
rect 9256 36928 9366 36988
rect 9256 36918 9366 36928
rect 10286 36928 10396 36988
rect 10286 36918 10396 36928
rect 13496 36998 13676 37478
rect 9776 36668 9886 36678
rect 9776 36608 9886 36668
rect 9966 36778 10236 36788
rect 9966 36628 10156 36778
rect 10156 36628 10236 36778
rect 9966 36618 10236 36628
rect 11956 36658 12156 36838
rect 14556 36618 14636 36838
rect 13976 36178 14256 36358
rect 14376 36158 14456 36378
rect 7446 36058 10656 36098
rect 7446 35988 7506 36058
rect 7506 35988 10606 36058
rect 10606 35988 10656 36058
rect 7446 35848 10656 35988
rect 12456 35838 12856 36018
rect 12976 35478 13356 35578
rect 12976 35418 13356 35478
rect 12216 35058 12396 35238
rect 13496 35058 13676 35238
rect 12536 34878 12576 34938
rect 12576 34878 12856 34938
rect 12536 34778 12856 34878
rect 17100 43820 17300 44000
rect 15780 43620 15960 43780
rect 16840 43420 16980 43540
rect 16100 43220 16240 43340
rect 12710 32886 12782 33214
rect 12556 32532 12876 32712
rect 5196 32192 5496 32372
rect 14576 32152 14656 32372
rect 7456 31332 10686 31492
rect 7456 31252 7466 31332
rect 7466 31252 10626 31332
rect 10626 31252 10686 31332
rect 7456 31222 10686 31252
rect 11616 31252 11836 31732
rect 13996 31712 14276 31892
rect 14396 31692 14476 31912
rect 7726 30742 7836 30752
rect 7726 30682 7836 30742
rect 7886 30852 8156 31062
rect 7886 30842 8106 30852
rect 8106 30842 8156 30852
rect 8246 31002 8356 31062
rect 8246 30992 8356 31002
rect 8756 30742 8866 30752
rect 8756 30682 8866 30742
rect 9276 31002 9386 31062
rect 9276 30992 9386 31002
rect 10306 31002 10416 31062
rect 10306 30992 10416 31002
rect 13516 31072 13696 31552
rect 9796 30742 9906 30752
rect 9796 30682 9906 30742
rect 9986 30852 10256 30862
rect 9986 30702 10176 30852
rect 10176 30702 10256 30852
rect 9986 30692 10256 30702
rect 11976 30732 12176 30912
rect 14576 30692 14656 30912
rect 13996 30252 14276 30432
rect 14396 30232 14476 30452
rect 7466 30132 10676 30172
rect 7466 30062 7526 30132
rect 7526 30062 10626 30132
rect 10626 30062 10676 30132
rect 7466 29922 10676 30062
rect 12476 29912 12876 30092
rect 12996 29552 13376 29652
rect 12996 29492 13376 29552
rect 11636 28992 11796 29272
rect 10856 28812 11796 28992
rect 12236 29132 12416 29312
rect 13516 29132 13696 29312
rect 12556 28952 12596 29012
rect 12596 28952 12876 29012
rect 12556 28852 12876 28952
rect 12824 26080 12898 26512
rect 12676 25828 12996 26008
rect 5316 25488 5616 25668
rect 14696 25448 14776 25668
rect 7576 24628 10806 24788
rect 7576 24548 7586 24628
rect 7586 24548 10746 24628
rect 10746 24548 10806 24628
rect 7576 24518 10806 24548
rect 11736 24548 11956 25028
rect 14116 25008 14396 25188
rect 14516 24988 14596 25208
rect 7846 24038 7956 24048
rect 7846 23978 7956 24038
rect 8006 24148 8276 24358
rect 8006 24138 8226 24148
rect 8226 24138 8276 24148
rect 8366 24298 8476 24358
rect 8366 24288 8476 24298
rect 8876 24038 8986 24048
rect 8876 23978 8986 24038
rect 9396 24298 9506 24358
rect 9396 24288 9506 24298
rect 10426 24298 10536 24358
rect 10426 24288 10536 24298
rect 13636 24368 13816 24848
rect 9916 24038 10026 24048
rect 9916 23978 10026 24038
rect 10106 24148 10376 24158
rect 10106 23998 10296 24148
rect 10296 23998 10376 24148
rect 10106 23988 10376 23998
rect 12096 24028 12296 24208
rect 14696 23988 14776 24208
rect 14116 23548 14396 23728
rect 14516 23528 14596 23748
rect 7586 23428 10796 23468
rect 7586 23358 7646 23428
rect 7646 23358 10746 23428
rect 10746 23358 10796 23428
rect 7586 23218 10796 23358
rect 12596 23208 12996 23388
rect 13116 22848 13496 22948
rect 13116 22788 13496 22848
rect 11756 22288 11916 22568
rect 10976 22108 11916 22288
rect 12356 22428 12536 22608
rect 13636 22428 13816 22608
rect 12676 22248 12716 22308
rect 12716 22248 12996 22308
rect 12676 22148 12996 22248
rect 16460 43000 16600 43140
rect 25432 38862 25502 39258
rect 25324 38576 25644 38756
rect 17964 38236 18264 38416
rect 27344 38196 27424 38416
rect 20224 37376 23454 37536
rect 20224 37296 20234 37376
rect 20234 37296 23394 37376
rect 23394 37296 23454 37376
rect 20224 37266 23454 37296
rect 24384 37296 24604 37776
rect 26764 37756 27044 37936
rect 27164 37736 27244 37956
rect 20494 36786 20604 36796
rect 20494 36726 20604 36786
rect 20654 36896 20924 37106
rect 20654 36886 20874 36896
rect 20874 36886 20924 36896
rect 21014 37046 21124 37106
rect 21014 37036 21124 37046
rect 21524 36786 21634 36796
rect 21524 36726 21634 36786
rect 22044 37046 22154 37106
rect 22044 37036 22154 37046
rect 23074 37046 23184 37106
rect 23074 37036 23184 37046
rect 26284 37116 26464 37596
rect 22564 36786 22674 36796
rect 22564 36726 22674 36786
rect 22754 36896 23024 36906
rect 22754 36746 22944 36896
rect 22944 36746 23024 36896
rect 22754 36736 23024 36746
rect 24744 36776 24944 36956
rect 27344 36736 27424 36956
rect 26764 36296 27044 36476
rect 27164 36276 27244 36496
rect 20234 36176 23444 36216
rect 20234 36106 20294 36176
rect 20294 36106 23394 36176
rect 23394 36106 23444 36176
rect 20234 35966 23444 36106
rect 25244 35956 25644 36136
rect 25764 35596 26144 35696
rect 25764 35536 26144 35596
rect 24404 35036 24564 35316
rect 23624 34856 24564 35036
rect 25004 35176 25184 35356
rect 26284 35176 26464 35356
rect 25324 34996 25364 35056
rect 25364 34996 25644 35056
rect 25324 34896 25644 34996
rect 25336 32804 25408 33132
rect 25288 32456 25608 32636
rect 17928 32116 18228 32296
rect 27308 32076 27388 32296
rect 20188 31256 23418 31416
rect 20188 31176 20198 31256
rect 20198 31176 23358 31256
rect 23358 31176 23418 31256
rect 20188 31146 23418 31176
rect 24348 31176 24568 31656
rect 26728 31636 27008 31816
rect 27128 31616 27208 31836
rect 20458 30666 20568 30676
rect 20458 30606 20568 30666
rect 20618 30776 20888 30986
rect 20618 30766 20838 30776
rect 20838 30766 20888 30776
rect 20978 30926 21088 30986
rect 20978 30916 21088 30926
rect 21488 30666 21598 30676
rect 21488 30606 21598 30666
rect 22008 30926 22118 30986
rect 22008 30916 22118 30926
rect 23038 30926 23148 30986
rect 23038 30916 23148 30926
rect 26248 30996 26428 31476
rect 22528 30666 22638 30676
rect 22528 30606 22638 30666
rect 22718 30776 22988 30786
rect 22718 30626 22908 30776
rect 22908 30626 22988 30776
rect 22718 30616 22988 30626
rect 24708 30656 24908 30836
rect 27308 30616 27388 30836
rect 26728 30176 27008 30356
rect 27128 30156 27208 30376
rect 20198 30056 23408 30096
rect 20198 29986 20258 30056
rect 20258 29986 23358 30056
rect 23358 29986 23408 30056
rect 20198 29846 23408 29986
rect 25208 29836 25608 30016
rect 25728 29476 26108 29576
rect 25728 29416 26108 29476
rect 24368 28916 24528 29196
rect 23588 28736 24528 28916
rect 24968 29056 25148 29236
rect 26248 29056 26428 29236
rect 25288 28876 25328 28936
rect 25328 28876 25608 28936
rect 25288 28776 25608 28876
rect 25518 25988 25586 26382
rect 25384 25698 25704 25878
rect 18024 25358 18324 25538
rect 27404 25318 27484 25538
rect 20284 24498 23514 24658
rect 20284 24418 20294 24498
rect 20294 24418 23454 24498
rect 23454 24418 23514 24498
rect 20284 24388 23514 24418
rect 24444 24418 24664 24898
rect 26824 24878 27104 25058
rect 27224 24858 27304 25078
rect 20554 23908 20664 23918
rect 20554 23848 20664 23908
rect 20714 24018 20984 24228
rect 20714 24008 20934 24018
rect 20934 24008 20984 24018
rect 21074 24168 21184 24228
rect 21074 24158 21184 24168
rect 21584 23908 21694 23918
rect 21584 23848 21694 23908
rect 22104 24168 22214 24228
rect 22104 24158 22214 24168
rect 23134 24168 23244 24228
rect 23134 24158 23244 24168
rect 26344 24238 26524 24718
rect 22624 23908 22734 23918
rect 22624 23848 22734 23908
rect 22814 24018 23084 24028
rect 22814 23868 23004 24018
rect 23004 23868 23084 24018
rect 22814 23858 23084 23868
rect 24804 23898 25004 24078
rect 27404 23858 27484 24078
rect 26824 23418 27104 23598
rect 27224 23398 27304 23618
rect 20294 23298 23504 23338
rect 20294 23228 20354 23298
rect 20354 23228 23454 23298
rect 23454 23228 23504 23298
rect 20294 23088 23504 23228
rect 25304 23078 25704 23258
rect 25824 22718 26204 22818
rect 25824 22658 26204 22718
rect 24464 22158 24624 22438
rect 23684 21978 24624 22158
rect 25064 22298 25244 22478
rect 26344 22298 26524 22478
rect 25384 22118 25424 22178
rect 25424 22118 25704 22178
rect 25384 22018 25704 22118
rect 12706 19126 12780 19464
rect 12552 18782 12872 18962
rect 25852 18942 25926 19334
rect 25734 18652 26054 18832
rect 5192 18442 5492 18622
rect 14572 18402 14652 18622
rect 18374 18312 18674 18492
rect 27754 18272 27834 18492
rect 7452 17582 10682 17742
rect 7452 17502 7462 17582
rect 7462 17502 10622 17582
rect 10622 17502 10682 17582
rect 7452 17472 10682 17502
rect 11612 17502 11832 17982
rect 13992 17962 14272 18142
rect 14392 17942 14472 18162
rect 7722 16992 7832 17002
rect 7722 16932 7832 16992
rect 7882 17102 8152 17312
rect 7882 17092 8102 17102
rect 8102 17092 8152 17102
rect 8242 17252 8352 17312
rect 8242 17242 8352 17252
rect 8752 16992 8862 17002
rect 8752 16932 8862 16992
rect 9272 17252 9382 17312
rect 9272 17242 9382 17252
rect 10302 17252 10412 17312
rect 10302 17242 10412 17252
rect 13512 17322 13692 17802
rect 20634 17452 23864 17612
rect 20634 17372 20644 17452
rect 20644 17372 23804 17452
rect 23804 17372 23864 17452
rect 20634 17342 23864 17372
rect 24794 17372 25014 17852
rect 27174 17832 27454 18012
rect 27574 17812 27654 18032
rect 9792 16992 9902 17002
rect 9792 16932 9902 16992
rect 9982 17102 10252 17112
rect 9982 16952 10172 17102
rect 10172 16952 10252 17102
rect 9982 16942 10252 16952
rect 11972 16982 12172 17162
rect 14572 16942 14652 17162
rect 20904 16862 21014 16872
rect 20904 16802 21014 16862
rect 21064 16972 21334 17182
rect 21064 16962 21284 16972
rect 21284 16962 21334 16972
rect 21424 17122 21534 17182
rect 21424 17112 21534 17122
rect 21934 16862 22044 16872
rect 21934 16802 22044 16862
rect 22454 17122 22564 17182
rect 22454 17112 22564 17122
rect 23484 17122 23594 17182
rect 23484 17112 23594 17122
rect 26694 17192 26874 17672
rect 22974 16862 23084 16872
rect 22974 16802 23084 16862
rect 23164 16972 23434 16982
rect 23164 16822 23354 16972
rect 23354 16822 23434 16972
rect 23164 16812 23434 16822
rect 25154 16852 25354 17032
rect 27754 16812 27834 17032
rect 13992 16502 14272 16682
rect 14392 16482 14472 16702
rect 7462 16382 10672 16422
rect 7462 16312 7522 16382
rect 7522 16312 10622 16382
rect 10622 16312 10672 16382
rect 7462 16172 10672 16312
rect 12472 16162 12872 16342
rect 27174 16372 27454 16552
rect 27574 16352 27654 16572
rect 20644 16252 23854 16292
rect 20644 16182 20704 16252
rect 20704 16182 23804 16252
rect 23804 16182 23854 16252
rect 20644 16042 23854 16182
rect 12992 15802 13372 15902
rect 12992 15742 13372 15802
rect 25654 16032 26054 16212
rect 11632 15242 11792 15522
rect 10852 15062 11792 15242
rect 12232 15382 12412 15562
rect 13512 15382 13692 15562
rect 12552 15202 12592 15262
rect 12592 15202 12872 15262
rect 12552 15102 12872 15202
rect 26174 15672 26554 15772
rect 26174 15612 26554 15672
rect 24814 15112 24974 15392
rect 24034 14932 24974 15112
rect 25414 15252 25594 15432
rect 26694 15252 26874 15432
rect 25734 15072 25774 15132
rect 25774 15072 26054 15132
rect 25734 14972 26054 15072
<< metal3 >>
rect 14960 44600 15140 44620
rect 14960 44480 14980 44600
rect 15120 44588 15140 44600
rect 29460 44600 29600 44620
rect 29460 44588 29480 44600
rect 15120 44495 29480 44588
rect 15120 44480 15140 44495
rect 14960 44460 15140 44480
rect 29460 44480 29480 44495
rect 29580 44480 29600 44600
rect 29460 44460 29600 44480
rect 17380 44400 17600 44420
rect 17380 44280 17400 44400
rect 17580 44386 17600 44400
rect 28720 44400 28880 44420
rect 28720 44386 28740 44400
rect 17580 44292 28740 44386
rect 17580 44280 17600 44292
rect 17380 44260 17600 44280
rect 28720 44280 28740 44292
rect 28860 44280 28880 44400
rect 28720 44260 28880 44280
rect 15380 44200 15600 44220
rect 15380 44040 15400 44200
rect 15580 44182 15600 44200
rect 27980 44200 28140 44220
rect 27980 44182 28000 44200
rect 15580 44088 28000 44182
rect 15580 44040 15600 44088
rect 15380 44020 15600 44040
rect 27980 44040 28000 44088
rect 28120 44040 28140 44200
rect 27980 44020 28140 44040
rect 17080 44000 17320 44020
rect 17080 43820 17100 44000
rect 17300 43956 17320 44000
rect 27220 44000 27420 44020
rect 27220 43956 27240 44000
rect 17300 43862 27240 43956
rect 17300 43820 17320 43862
rect 17080 43800 17320 43820
rect 27220 43820 27240 43862
rect 27400 43820 27420 44000
rect 27220 43800 27420 43820
rect 15760 43780 15980 43800
rect 15760 43620 15780 43780
rect 15960 43728 15980 43780
rect 26500 43760 26680 43780
rect 26500 43728 26520 43760
rect 15960 43634 26520 43728
rect 15960 43620 15980 43634
rect 15760 43600 15980 43620
rect 26500 43620 26520 43634
rect 26660 43620 26680 43760
rect 26500 43600 26680 43620
rect 16820 43540 17000 43560
rect 16820 43420 16840 43540
rect 16980 43524 17000 43540
rect 25720 43540 25960 43560
rect 25720 43524 25760 43540
rect 16980 43430 25760 43524
rect 16980 43420 17000 43430
rect 16820 43400 17000 43420
rect 25720 43420 25760 43430
rect 25940 43420 25960 43540
rect 25720 43400 25960 43420
rect 16080 43340 16260 43360
rect 16080 43220 16100 43340
rect 16240 43320 16260 43340
rect 25000 43340 25220 43360
rect 25000 43320 25020 43340
rect 16240 43226 25020 43320
rect 16240 43220 16260 43226
rect 16080 43200 16260 43220
rect 25000 43220 25020 43226
rect 25200 43220 25220 43340
rect 25000 43200 25220 43220
rect 16440 43140 16620 43160
rect 16440 43000 16460 43140
rect 16600 43128 16620 43140
rect 24260 43140 24480 43160
rect 24260 43128 24280 43140
rect 16600 43034 24280 43128
rect 16600 43000 16620 43034
rect 16440 42980 16620 43000
rect 24260 43000 24280 43034
rect 24460 43000 24480 43140
rect 24260 42980 24480 43000
rect 25304 39258 25664 39276
rect 12516 39108 12876 39158
rect 13956 39120 14276 39158
rect 17944 39120 18284 39136
rect 5156 39012 5496 39018
rect 2490 38596 5496 39012
rect 2490 2600 2906 38596
rect 5156 38298 5496 38596
rect 5156 38118 5176 38298
rect 5476 38118 5496 38298
rect 5156 37058 5496 38118
rect 12516 38710 12656 39108
rect 12734 38710 12876 39108
rect 13930 38800 18284 39120
rect 12516 38638 12876 38710
rect 12516 38458 12536 38638
rect 12856 38458 12876 38638
rect 5616 37938 11316 37998
rect 5616 37198 5676 37938
rect 11236 37198 11316 37938
rect 5616 37148 7436 37198
rect 10666 37148 11316 37198
rect 5616 37138 11316 37148
rect 11576 37658 11836 37678
rect 11576 37178 11596 37658
rect 11816 37178 11836 37658
rect 11576 37118 11836 37178
rect 5156 36988 8146 37058
rect 11576 37018 12176 37118
rect 10036 36998 12176 37018
rect 5156 36768 7866 36988
rect 8136 36768 8146 36988
rect 5156 36758 8146 36768
rect 7476 36748 8146 36758
rect 8206 36988 12176 36998
rect 8206 36918 8226 36988
rect 8336 36918 9256 36988
rect 9366 36918 10286 36988
rect 10396 36918 12176 36988
rect 8206 36908 10702 36918
rect 8206 36748 9866 36908
rect 10282 36848 10702 36908
rect 9956 36788 10702 36848
rect 7696 36678 9896 36688
rect 7696 36608 7706 36678
rect 7816 36608 8736 36678
rect 8846 36608 9776 36678
rect 9886 36608 9896 36678
rect 7696 36598 9896 36608
rect 8236 36438 9896 36598
rect 9956 36618 9966 36788
rect 10236 36618 10702 36788
rect 11936 36838 12176 36918
rect 11936 36658 11956 36838
rect 12156 36658 12176 36838
rect 11936 36638 12176 36658
rect 9956 36474 10702 36618
rect 9956 36458 10626 36474
rect 5616 36098 11316 36128
rect 5616 36078 7446 36098
rect 10656 36078 11316 36098
rect 12516 36078 12876 38458
rect 5616 35258 5676 36078
rect 11256 35258 11316 36078
rect 5616 35198 11316 35258
rect 12196 36018 12876 36078
rect 12196 35838 12456 36018
rect 12856 35838 12876 36018
rect 12196 35758 12876 35838
rect 12956 37978 13376 37998
rect 12956 37158 12976 37978
rect 13356 37158 13376 37978
rect 13956 37818 14276 38800
rect 17944 38416 18284 38800
rect 14536 38298 14656 38318
rect 14536 38078 14556 38298
rect 14636 38078 14656 38298
rect 14536 37978 14656 38078
rect 13956 37638 13976 37818
rect 14256 37638 14276 37818
rect 12196 35238 12416 35758
rect 12196 35058 12216 35238
rect 12396 35058 12416 35238
rect 12196 35038 12416 35058
rect 12516 35578 12876 35598
rect 12516 35218 12536 35578
rect 12856 35218 12876 35578
rect 12956 35578 13376 37158
rect 12956 35418 12976 35578
rect 13356 35418 13376 35578
rect 12956 35398 13376 35418
rect 13476 37478 13696 37498
rect 13476 36998 13496 37478
rect 13676 36998 13696 37478
rect 12516 34938 12876 35218
rect 13476 35238 13696 36998
rect 13956 36358 14276 37638
rect 13956 36178 13976 36358
rect 14256 36178 14276 36358
rect 13956 36158 14276 36178
rect 14356 37838 14476 37858
rect 14356 37618 14376 37838
rect 14456 37618 14476 37838
rect 14356 36378 14476 37618
rect 14536 37158 14556 37978
rect 14636 37158 14656 37978
rect 14536 36838 14656 37158
rect 17944 38236 17964 38416
rect 18264 38236 18284 38416
rect 17944 37176 18284 38236
rect 25304 38862 25432 39258
rect 25502 38862 25664 39258
rect 25304 38756 25664 38862
rect 25304 38576 25324 38756
rect 25644 38576 25664 38756
rect 18404 38056 24104 38116
rect 18404 37316 18464 38056
rect 24024 37316 24104 38056
rect 18404 37266 20224 37316
rect 23454 37266 24104 37316
rect 18404 37256 24104 37266
rect 24364 37776 24624 37796
rect 24364 37296 24384 37776
rect 24604 37296 24624 37776
rect 24364 37236 24624 37296
rect 17944 37106 20934 37176
rect 24364 37136 24964 37236
rect 22824 37116 24964 37136
rect 17944 36886 20654 37106
rect 20924 36886 20934 37106
rect 17944 36876 20934 36886
rect 20264 36866 20934 36876
rect 20994 37106 24964 37116
rect 20994 37036 21014 37106
rect 21124 37036 22044 37106
rect 22154 37036 23074 37106
rect 23184 37036 24964 37106
rect 20994 37026 23194 37036
rect 20994 36866 22654 37026
rect 22744 36956 23414 36966
rect 24724 36956 24964 37036
rect 22744 36906 24584 36956
rect 14536 36618 14556 36838
rect 14636 36618 14656 36838
rect 20484 36796 22684 36806
rect 20484 36726 20494 36796
rect 20604 36726 21524 36796
rect 21634 36726 22564 36796
rect 22674 36726 22684 36796
rect 20484 36716 22684 36726
rect 14536 36598 14656 36618
rect 21024 36556 22684 36716
rect 22744 36736 22754 36906
rect 23024 36736 24584 36906
rect 24724 36776 24744 36956
rect 24944 36776 24964 36956
rect 24724 36756 24964 36776
rect 22744 36576 24584 36736
rect 14356 36158 14376 36378
rect 14456 36158 14476 36378
rect 13476 35058 13496 35238
rect 13676 35058 13696 35238
rect 14356 36118 14476 36158
rect 14356 35218 14376 36118
rect 14456 35218 14476 36118
rect 18404 36216 24104 36246
rect 18404 36196 20234 36216
rect 23444 36196 24104 36216
rect 18404 35376 18464 36196
rect 24044 35376 24104 36196
rect 18404 35316 24104 35376
rect 24384 35316 24584 36576
rect 25304 36196 25664 38576
rect 26744 39269 27064 39276
rect 29335 39269 29658 39272
rect 26744 38951 29658 39269
rect 14356 35198 14476 35218
rect 13476 35038 13696 35058
rect 24384 35056 24404 35316
rect 12516 34778 12536 34938
rect 12856 34778 12876 34938
rect 23604 35036 24404 35056
rect 23604 34856 23624 35036
rect 24564 34856 24584 35316
rect 24984 36136 25664 36196
rect 24984 35956 25244 36136
rect 25644 35956 25664 36136
rect 24984 35876 25664 35956
rect 25744 38096 26164 38116
rect 25744 37276 25764 38096
rect 26144 37276 26164 38096
rect 26744 37936 27064 38951
rect 27324 38416 27444 38436
rect 27324 38196 27344 38416
rect 27424 38196 27444 38416
rect 27324 38096 27444 38196
rect 26744 37756 26764 37936
rect 27044 37756 27064 37936
rect 24984 35356 25204 35876
rect 24984 35176 25004 35356
rect 25184 35176 25204 35356
rect 24984 35156 25204 35176
rect 25304 35696 25664 35716
rect 25304 35336 25324 35696
rect 25644 35336 25664 35696
rect 25744 35696 26164 37276
rect 25744 35536 25764 35696
rect 26144 35536 26164 35696
rect 25744 35516 26164 35536
rect 26264 37596 26484 37616
rect 26264 37116 26284 37596
rect 26464 37116 26484 37596
rect 25304 35056 25664 35336
rect 26264 35356 26484 37116
rect 26744 36476 27064 37756
rect 26744 36296 26764 36476
rect 27044 36296 27064 36476
rect 26744 36276 27064 36296
rect 27144 37956 27264 37976
rect 27144 37736 27164 37956
rect 27244 37736 27264 37956
rect 27144 36496 27264 37736
rect 27324 37276 27344 38096
rect 27424 37276 27444 38096
rect 27324 36956 27444 37276
rect 27324 36736 27344 36956
rect 27424 36736 27444 36956
rect 27324 36716 27444 36736
rect 27144 36276 27164 36496
rect 27244 36276 27264 36496
rect 26264 35176 26284 35356
rect 26464 35176 26484 35356
rect 27144 36236 27264 36276
rect 27144 35336 27164 36236
rect 27244 35336 27264 36236
rect 27144 35316 27264 35336
rect 26264 35156 26484 35176
rect 25304 34896 25324 35056
rect 25644 34896 25664 35056
rect 25304 34876 25664 34896
rect 23604 34836 24584 34856
rect 12516 34758 12876 34778
rect 29335 34518 29658 38951
rect 5090 34198 29658 34518
rect 5092 32668 5519 34198
rect 29335 34197 29658 34198
rect 12536 33214 12896 33232
rect 12536 32886 12710 33214
rect 12782 32886 12896 33214
rect 12536 32712 12896 32886
rect 5094 32372 5516 32668
rect 5094 32368 5196 32372
rect 5176 32192 5196 32368
rect 5496 32192 5516 32372
rect 5176 31132 5516 32192
rect 12536 32532 12556 32712
rect 12876 32532 12896 32712
rect 5636 32012 11336 32072
rect 5636 31272 5696 32012
rect 11256 31272 11336 32012
rect 5636 31222 7456 31272
rect 10686 31222 11336 31272
rect 5636 31212 11336 31222
rect 11596 31732 11856 31752
rect 11596 31252 11616 31732
rect 11836 31252 11856 31732
rect 11596 31192 11856 31252
rect 5176 31062 8166 31132
rect 11596 31092 12196 31192
rect 10056 31072 12196 31092
rect 5176 30842 7886 31062
rect 8156 30842 8166 31062
rect 5176 30832 8166 30842
rect 7496 30822 8166 30832
rect 8226 31062 12196 31072
rect 8226 30992 8246 31062
rect 8356 30992 9276 31062
rect 9386 30992 10306 31062
rect 10416 30992 12196 31062
rect 8226 30982 10426 30992
rect 8226 30822 9886 30982
rect 9976 30912 10646 30922
rect 11956 30912 12196 30992
rect 9976 30862 11816 30912
rect 7716 30752 9916 30762
rect 7716 30682 7726 30752
rect 7836 30682 8756 30752
rect 8866 30682 9796 30752
rect 9906 30682 9916 30752
rect 7716 30672 9916 30682
rect 8256 30512 9916 30672
rect 9976 30692 9986 30862
rect 10256 30692 11816 30862
rect 11956 30732 11976 30912
rect 12176 30732 12196 30912
rect 11956 30712 12196 30732
rect 9976 30532 11816 30692
rect 5636 30172 11336 30202
rect 5636 30152 7466 30172
rect 10676 30152 11336 30172
rect 5636 29332 5696 30152
rect 11276 29332 11336 30152
rect 5636 29272 11336 29332
rect 11616 29272 11816 30532
rect 12536 30152 12896 32532
rect 13976 32994 14296 33232
rect 25268 33132 25628 33156
rect 17908 32994 18248 33016
rect 13976 32654 18248 32994
rect 11616 29012 11636 29272
rect 10836 28992 11636 29012
rect 10836 28812 10856 28992
rect 11796 28812 11816 29272
rect 12216 30092 12896 30152
rect 12216 29912 12476 30092
rect 12876 29912 12896 30092
rect 12216 29832 12896 29912
rect 12976 32052 13396 32072
rect 12976 31232 12996 32052
rect 13376 31232 13396 32052
rect 13976 31892 14296 32654
rect 14556 32372 14676 32392
rect 14556 32152 14576 32372
rect 14656 32152 14676 32372
rect 14556 32052 14676 32152
rect 13976 31712 13996 31892
rect 14276 31712 14296 31892
rect 12216 29312 12436 29832
rect 12216 29132 12236 29312
rect 12416 29132 12436 29312
rect 12216 29112 12436 29132
rect 12536 29652 12896 29672
rect 12536 29292 12556 29652
rect 12876 29292 12896 29652
rect 12976 29652 13396 31232
rect 12976 29492 12996 29652
rect 13376 29492 13396 29652
rect 12976 29472 13396 29492
rect 13496 31552 13716 31572
rect 13496 31072 13516 31552
rect 13696 31072 13716 31552
rect 12536 29012 12896 29292
rect 13496 29312 13716 31072
rect 13976 30432 14296 31712
rect 13976 30252 13996 30432
rect 14276 30252 14296 30432
rect 13976 30232 14296 30252
rect 14376 31912 14496 31932
rect 14376 31692 14396 31912
rect 14476 31692 14496 31912
rect 14376 30452 14496 31692
rect 14556 31232 14576 32052
rect 14656 31232 14676 32052
rect 14556 30912 14676 31232
rect 14556 30692 14576 30912
rect 14656 30692 14676 30912
rect 17908 32296 18248 32654
rect 17908 32116 17928 32296
rect 18228 32116 18248 32296
rect 17908 31056 18248 32116
rect 25268 32804 25336 33132
rect 25408 32804 25628 33132
rect 25268 32636 25628 32804
rect 25268 32456 25288 32636
rect 25608 32456 25628 32636
rect 18368 31936 24068 31996
rect 18368 31196 18428 31936
rect 23988 31196 24068 31936
rect 18368 31146 20188 31196
rect 23418 31146 24068 31196
rect 18368 31136 24068 31146
rect 24328 31656 24588 31676
rect 24328 31176 24348 31656
rect 24568 31176 24588 31656
rect 24328 31116 24588 31176
rect 17908 30986 20898 31056
rect 24328 31016 24928 31116
rect 22788 30996 24928 31016
rect 17908 30766 20618 30986
rect 20888 30766 20898 30986
rect 17908 30756 20898 30766
rect 20228 30746 20898 30756
rect 20958 30986 24928 30996
rect 20958 30916 20978 30986
rect 21088 30916 22008 30986
rect 22118 30916 23038 30986
rect 23148 30916 24928 30986
rect 20958 30906 23158 30916
rect 20958 30746 22618 30906
rect 22708 30836 23378 30846
rect 24688 30836 24928 30916
rect 22708 30786 24548 30836
rect 14556 30672 14676 30692
rect 20448 30676 22648 30686
rect 20448 30606 20458 30676
rect 20568 30606 21488 30676
rect 21598 30606 22528 30676
rect 22638 30606 22648 30676
rect 20448 30596 22648 30606
rect 14376 30232 14396 30452
rect 14476 30232 14496 30452
rect 20988 30436 22648 30596
rect 22708 30616 22718 30786
rect 22988 30616 24548 30786
rect 24688 30656 24708 30836
rect 24908 30656 24928 30836
rect 24688 30636 24928 30656
rect 22708 30456 24548 30616
rect 13496 29132 13516 29312
rect 13696 29132 13716 29312
rect 14376 30192 14496 30232
rect 14376 29292 14396 30192
rect 14476 29292 14496 30192
rect 14376 29272 14496 29292
rect 18368 30096 24068 30126
rect 18368 30076 20198 30096
rect 23408 30076 24068 30096
rect 18368 29256 18428 30076
rect 24008 29256 24068 30076
rect 18368 29196 24068 29256
rect 24348 29196 24548 30456
rect 25268 30076 25628 32456
rect 26708 32836 29522 33156
rect 13496 29112 13716 29132
rect 12536 28852 12556 29012
rect 12876 28852 12896 29012
rect 24348 28936 24368 29196
rect 12536 28832 12896 28852
rect 23568 28916 24368 28936
rect 10836 28792 11816 28812
rect 23568 28736 23588 28916
rect 24528 28736 24548 29196
rect 24948 30016 25628 30076
rect 24948 29836 25208 30016
rect 25608 29836 25628 30016
rect 24948 29756 25628 29836
rect 25708 31976 26128 31996
rect 25708 31156 25728 31976
rect 26108 31156 26128 31976
rect 26708 31816 27028 32836
rect 27288 32296 27408 32316
rect 27288 32076 27308 32296
rect 27388 32076 27408 32296
rect 27288 31976 27408 32076
rect 26708 31636 26728 31816
rect 27008 31636 27028 31816
rect 24948 29236 25168 29756
rect 24948 29056 24968 29236
rect 25148 29056 25168 29236
rect 24948 29036 25168 29056
rect 25268 29576 25628 29596
rect 25268 29216 25288 29576
rect 25608 29216 25628 29576
rect 25708 29576 26128 31156
rect 25708 29416 25728 29576
rect 26108 29416 26128 29576
rect 25708 29396 26128 29416
rect 26228 31476 26448 31496
rect 26228 30996 26248 31476
rect 26428 30996 26448 31476
rect 25268 28936 25628 29216
rect 26228 29236 26448 30996
rect 26708 30356 27028 31636
rect 26708 30176 26728 30356
rect 27008 30176 27028 30356
rect 26708 30156 27028 30176
rect 27108 31836 27228 31856
rect 27108 31616 27128 31836
rect 27208 31616 27228 31836
rect 27108 30376 27228 31616
rect 27288 31156 27308 31976
rect 27388 31156 27408 31976
rect 27288 30836 27408 31156
rect 27288 30616 27308 30836
rect 27388 30616 27408 30836
rect 27288 30596 27408 30616
rect 27108 30156 27128 30376
rect 27208 30156 27228 30376
rect 26228 29056 26248 29236
rect 26428 29056 26448 29236
rect 27108 30116 27228 30156
rect 27108 29216 27128 30116
rect 27208 29216 27228 30116
rect 27108 29196 27228 29216
rect 26228 29036 26448 29056
rect 25268 28776 25288 28936
rect 25608 28776 25628 28936
rect 25268 28756 25628 28776
rect 23568 28716 24548 28736
rect 29204 28398 29520 32836
rect 5290 28082 29520 28398
rect 5296 25668 5636 28082
rect 5296 25488 5316 25668
rect 5616 25488 5636 25668
rect 5296 24428 5636 25488
rect 12656 26512 13016 26528
rect 12656 26080 12824 26512
rect 12898 26080 13016 26512
rect 12656 26008 13016 26080
rect 12656 25828 12676 26008
rect 12996 25828 13016 26008
rect 5756 25308 11456 25368
rect 5756 24568 5816 25308
rect 11376 24568 11456 25308
rect 5756 24518 7576 24568
rect 10806 24518 11456 24568
rect 5756 24508 11456 24518
rect 11716 25028 11976 25048
rect 11716 24548 11736 25028
rect 11956 24548 11976 25028
rect 11716 24488 11976 24548
rect 5296 24358 8286 24428
rect 11716 24388 12316 24488
rect 10176 24368 12316 24388
rect 5296 24138 8006 24358
rect 8276 24138 8286 24358
rect 5296 24128 8286 24138
rect 7616 24118 8286 24128
rect 8346 24358 12316 24368
rect 8346 24288 8366 24358
rect 8476 24288 9396 24358
rect 9506 24288 10426 24358
rect 10536 24288 12316 24358
rect 8346 24278 10546 24288
rect 8346 24118 10006 24278
rect 10096 24208 10766 24218
rect 12076 24208 12316 24288
rect 10096 24158 11936 24208
rect 7836 24048 10036 24058
rect 7836 23978 7846 24048
rect 7956 23978 8876 24048
rect 8986 23978 9916 24048
rect 10026 23978 10036 24048
rect 7836 23968 10036 23978
rect 8376 23808 10036 23968
rect 10096 23988 10106 24158
rect 10376 23988 11936 24158
rect 12076 24028 12096 24208
rect 12296 24028 12316 24208
rect 12076 24008 12316 24028
rect 10096 23828 11936 23988
rect 5756 23468 11456 23498
rect 5756 23448 7586 23468
rect 10796 23448 11456 23468
rect 5756 22628 5816 23448
rect 11396 22628 11456 23448
rect 5756 22568 11456 22628
rect 11736 22568 11936 23828
rect 12656 23448 13016 25828
rect 14096 26280 14416 26528
rect 25364 26382 25724 26398
rect 14096 25960 18366 26280
rect 25364 25988 25518 26382
rect 25586 25988 25724 26382
rect 11736 22308 11756 22568
rect 10956 22288 11756 22308
rect 10956 22108 10976 22288
rect 11916 22108 11936 22568
rect 12336 23388 13016 23448
rect 12336 23208 12596 23388
rect 12996 23208 13016 23388
rect 12336 23128 13016 23208
rect 13096 25348 13516 25368
rect 13096 24528 13116 25348
rect 13496 24528 13516 25348
rect 14096 25188 14416 25960
rect 14676 25668 14796 25688
rect 14676 25448 14696 25668
rect 14776 25448 14796 25668
rect 14676 25348 14796 25448
rect 14096 25008 14116 25188
rect 14396 25008 14416 25188
rect 12336 22608 12556 23128
rect 12336 22428 12356 22608
rect 12536 22428 12556 22608
rect 12336 22408 12556 22428
rect 12656 22948 13016 22968
rect 12656 22588 12676 22948
rect 12996 22588 13016 22948
rect 13096 22948 13516 24528
rect 13096 22788 13116 22948
rect 13496 22788 13516 22948
rect 13096 22768 13516 22788
rect 13616 24848 13836 24868
rect 13616 24368 13636 24848
rect 13816 24368 13836 24848
rect 12656 22308 13016 22588
rect 13616 22608 13836 24368
rect 14096 23728 14416 25008
rect 14096 23548 14116 23728
rect 14396 23548 14416 23728
rect 14096 23528 14416 23548
rect 14496 25208 14616 25228
rect 14496 24988 14516 25208
rect 14596 24988 14616 25208
rect 14496 23748 14616 24988
rect 14676 24528 14696 25348
rect 14776 24528 14796 25348
rect 14676 24208 14796 24528
rect 14676 23988 14696 24208
rect 14776 23988 14796 24208
rect 18004 25538 18344 25960
rect 18004 25358 18024 25538
rect 18324 25358 18344 25538
rect 18004 24298 18344 25358
rect 25364 25878 25724 25988
rect 25364 25698 25384 25878
rect 25704 25698 25724 25878
rect 18464 25178 24164 25238
rect 18464 24438 18524 25178
rect 24084 24438 24164 25178
rect 18464 24388 20284 24438
rect 23514 24388 24164 24438
rect 18464 24378 24164 24388
rect 24424 24898 24684 24918
rect 24424 24418 24444 24898
rect 24664 24418 24684 24898
rect 24424 24358 24684 24418
rect 18004 24228 20994 24298
rect 24424 24258 25024 24358
rect 22884 24238 25024 24258
rect 18004 24008 20714 24228
rect 20984 24008 20994 24228
rect 18004 23998 20994 24008
rect 20324 23988 20994 23998
rect 21054 24228 25024 24238
rect 21054 24158 21074 24228
rect 21184 24158 22104 24228
rect 22214 24158 23134 24228
rect 23244 24158 25024 24228
rect 21054 24148 23254 24158
rect 21054 23988 22714 24148
rect 22804 24078 23474 24088
rect 24784 24078 25024 24158
rect 22804 24028 24644 24078
rect 14676 23968 14796 23988
rect 20544 23918 22744 23928
rect 20544 23848 20554 23918
rect 20664 23848 21584 23918
rect 21694 23848 22624 23918
rect 22734 23848 22744 23918
rect 20544 23838 22744 23848
rect 14496 23528 14516 23748
rect 14596 23528 14616 23748
rect 21084 23678 22744 23838
rect 22804 23858 22814 24028
rect 23084 23858 24644 24028
rect 24784 23898 24804 24078
rect 25004 23898 25024 24078
rect 24784 23878 25024 23898
rect 22804 23698 24644 23858
rect 13616 22428 13636 22608
rect 13816 22428 13836 22608
rect 14496 23488 14616 23528
rect 14496 22588 14516 23488
rect 14596 22588 14616 23488
rect 14496 22568 14616 22588
rect 18464 23338 24164 23368
rect 18464 23318 20294 23338
rect 23504 23318 24164 23338
rect 18464 22498 18524 23318
rect 24104 22498 24164 23318
rect 18464 22438 24164 22498
rect 24444 22438 24644 23698
rect 25364 23318 25724 25698
rect 26804 26266 27124 26398
rect 26804 25946 29360 26266
rect 13616 22408 13836 22428
rect 12656 22148 12676 22308
rect 12996 22148 13016 22308
rect 24444 22178 24464 22438
rect 12656 22128 13016 22148
rect 23664 22158 24464 22178
rect 10956 22088 11936 22108
rect 23664 21978 23684 22158
rect 24624 21978 24644 22438
rect 25044 23258 25724 23318
rect 25044 23078 25304 23258
rect 25704 23078 25724 23258
rect 25044 22998 25724 23078
rect 25804 25218 26224 25238
rect 25804 24398 25824 25218
rect 26204 24398 26224 25218
rect 26804 25058 27124 25946
rect 27384 25538 27504 25558
rect 27384 25318 27404 25538
rect 27484 25318 27504 25538
rect 27384 25218 27504 25318
rect 26804 24878 26824 25058
rect 27104 24878 27124 25058
rect 25044 22478 25264 22998
rect 25044 22298 25064 22478
rect 25244 22298 25264 22478
rect 25044 22278 25264 22298
rect 25364 22818 25724 22838
rect 25364 22458 25384 22818
rect 25704 22458 25724 22818
rect 25804 22818 26224 24398
rect 25804 22658 25824 22818
rect 26204 22658 26224 22818
rect 25804 22638 26224 22658
rect 26324 24718 26544 24738
rect 26324 24238 26344 24718
rect 26524 24238 26544 24718
rect 25364 22178 25724 22458
rect 26324 22478 26544 24238
rect 26804 23598 27124 24878
rect 26804 23418 26824 23598
rect 27104 23418 27124 23598
rect 26804 23398 27124 23418
rect 27204 25078 27324 25098
rect 27204 24858 27224 25078
rect 27304 24858 27324 25078
rect 27204 23618 27324 24858
rect 27384 24398 27404 25218
rect 27484 24398 27504 25218
rect 27384 24078 27504 24398
rect 27384 23858 27404 24078
rect 27484 23858 27504 24078
rect 27384 23838 27504 23858
rect 27204 23398 27224 23618
rect 27304 23398 27324 23618
rect 26324 22298 26344 22478
rect 26524 22298 26544 22478
rect 27204 23358 27324 23398
rect 27204 22458 27224 23358
rect 27304 22458 27324 23358
rect 27204 22438 27324 22458
rect 26324 22278 26544 22298
rect 25364 22018 25384 22178
rect 25704 22018 25724 22178
rect 25364 21998 25724 22018
rect 23664 21958 24644 21978
rect 5172 21674 5512 21690
rect 29040 21674 29360 25946
rect 5172 21354 29360 21674
rect 5172 18622 5512 21354
rect 5172 18442 5192 18622
rect 5492 18442 5512 18622
rect 5172 17382 5512 18442
rect 12532 19464 12892 19482
rect 12532 19126 12706 19464
rect 12780 19126 12892 19464
rect 12532 18962 12892 19126
rect 12532 18782 12552 18962
rect 12872 18782 12892 18962
rect 5632 18262 11332 18322
rect 5632 17522 5692 18262
rect 11252 17522 11332 18262
rect 5632 17472 7452 17522
rect 10682 17472 11332 17522
rect 5632 17462 11332 17472
rect 11592 17982 11852 18002
rect 11592 17502 11612 17982
rect 11832 17502 11852 17982
rect 11592 17442 11852 17502
rect 5172 17312 8162 17382
rect 11592 17342 12192 17442
rect 10052 17322 12192 17342
rect 5172 17092 7882 17312
rect 8152 17092 8162 17312
rect 5172 17082 8162 17092
rect 7492 17072 8162 17082
rect 8222 17312 12192 17322
rect 8222 17242 8242 17312
rect 8352 17242 9272 17312
rect 9382 17242 10302 17312
rect 10412 17242 12192 17312
rect 8222 17232 10422 17242
rect 8222 17072 9882 17232
rect 9972 17162 10642 17172
rect 11952 17162 12192 17242
rect 9972 17112 11812 17162
rect 7712 17002 9912 17012
rect 7712 16932 7722 17002
rect 7832 16932 8752 17002
rect 8862 16932 9792 17002
rect 9902 16932 9912 17002
rect 7712 16922 9912 16932
rect 8252 16762 9912 16922
rect 9972 16942 9982 17112
rect 10252 16942 11812 17112
rect 11952 16982 11972 17162
rect 12172 16982 12192 17162
rect 11952 16962 12192 16982
rect 9972 16782 11812 16942
rect 5632 16422 11332 16452
rect 5632 16402 7462 16422
rect 10672 16402 11332 16422
rect 5632 15582 5692 16402
rect 11272 15582 11332 16402
rect 5632 15522 11332 15582
rect 11612 15522 11812 16782
rect 12532 16402 12892 18782
rect 13972 19456 14292 19482
rect 13972 19212 18688 19456
rect 25714 19334 26074 19352
rect 13972 19136 18694 19212
rect 11612 15262 11632 15522
rect 10832 15242 11632 15262
rect 10832 15062 10852 15242
rect 11792 15062 11812 15522
rect 12212 16342 12892 16402
rect 12212 16162 12472 16342
rect 12872 16162 12892 16342
rect 12212 16082 12892 16162
rect 12972 18302 13392 18322
rect 12972 17482 12992 18302
rect 13372 17482 13392 18302
rect 13972 18142 14292 19136
rect 14552 18622 14672 18642
rect 14552 18402 14572 18622
rect 14652 18402 14672 18622
rect 14552 18302 14672 18402
rect 13972 17962 13992 18142
rect 14272 17962 14292 18142
rect 12212 15562 12432 16082
rect 12212 15382 12232 15562
rect 12412 15382 12432 15562
rect 12212 15362 12432 15382
rect 12532 15902 12892 15922
rect 12532 15542 12552 15902
rect 12872 15542 12892 15902
rect 12972 15902 13392 17482
rect 12972 15742 12992 15902
rect 13372 15742 13392 15902
rect 12972 15722 13392 15742
rect 13492 17802 13712 17822
rect 13492 17322 13512 17802
rect 13692 17322 13712 17802
rect 12532 15262 12892 15542
rect 13492 15562 13712 17322
rect 13972 16682 14292 17962
rect 13972 16502 13992 16682
rect 14272 16502 14292 16682
rect 13972 16482 14292 16502
rect 14372 18162 14492 18182
rect 14372 17942 14392 18162
rect 14472 17942 14492 18162
rect 14372 16702 14492 17942
rect 14552 17482 14572 18302
rect 14652 17482 14672 18302
rect 14552 17162 14672 17482
rect 14552 16942 14572 17162
rect 14652 16942 14672 17162
rect 18354 18492 18694 19136
rect 18354 18312 18374 18492
rect 18674 18312 18694 18492
rect 18354 17252 18694 18312
rect 25714 18942 25852 19334
rect 25926 18942 26074 19334
rect 25714 18832 26074 18942
rect 25714 18652 25734 18832
rect 26054 18652 26074 18832
rect 18814 18132 24514 18192
rect 18814 17392 18874 18132
rect 24434 17392 24514 18132
rect 18814 17342 20634 17392
rect 23864 17342 24514 17392
rect 18814 17332 24514 17342
rect 24774 17852 25034 17872
rect 24774 17372 24794 17852
rect 25014 17372 25034 17852
rect 24774 17312 25034 17372
rect 18354 17182 21344 17252
rect 24774 17212 25374 17312
rect 23234 17192 25374 17212
rect 18354 16962 21064 17182
rect 21334 16962 21344 17182
rect 18354 16952 21344 16962
rect 20674 16942 21344 16952
rect 21404 17182 25374 17192
rect 21404 17112 21424 17182
rect 21534 17112 22454 17182
rect 22564 17112 23484 17182
rect 23594 17112 25374 17182
rect 21404 17102 23604 17112
rect 21404 16942 23064 17102
rect 23154 17032 23824 17042
rect 25134 17032 25374 17112
rect 23154 16982 24994 17032
rect 14552 16922 14672 16942
rect 20894 16872 23094 16882
rect 20894 16802 20904 16872
rect 21014 16802 21934 16872
rect 22044 16802 22974 16872
rect 23084 16802 23094 16872
rect 20894 16792 23094 16802
rect 14372 16482 14392 16702
rect 14472 16482 14492 16702
rect 21434 16632 23094 16792
rect 23154 16812 23164 16982
rect 23434 16812 24994 16982
rect 25134 16852 25154 17032
rect 25354 16852 25374 17032
rect 25134 16832 25374 16852
rect 23154 16652 24994 16812
rect 13492 15382 13512 15562
rect 13692 15382 13712 15562
rect 14372 16442 14492 16482
rect 14372 15542 14392 16442
rect 14472 15542 14492 16442
rect 14372 15522 14492 15542
rect 18814 16292 24514 16322
rect 18814 16272 20644 16292
rect 23854 16272 24514 16292
rect 18814 15452 18874 16272
rect 24454 15452 24514 16272
rect 18814 15392 24514 15452
rect 24794 15392 24994 16652
rect 25714 16272 26074 18652
rect 27154 19032 29640 19352
rect 13492 15362 13712 15382
rect 12532 15102 12552 15262
rect 12872 15102 12892 15262
rect 24794 15132 24814 15392
rect 12532 15082 12892 15102
rect 24014 15112 24814 15132
rect 10832 15042 11812 15062
rect 24014 14932 24034 15112
rect 24974 14932 24994 15392
rect 25394 16212 26074 16272
rect 25394 16032 25654 16212
rect 26054 16032 26074 16212
rect 25394 15952 26074 16032
rect 26154 18172 26574 18192
rect 26154 17352 26174 18172
rect 26554 17352 26574 18172
rect 27154 18012 27474 19032
rect 27734 18492 27854 18512
rect 27734 18272 27754 18492
rect 27834 18272 27854 18492
rect 27734 18172 27854 18272
rect 27154 17832 27174 18012
rect 27454 17832 27474 18012
rect 25394 15432 25614 15952
rect 25394 15252 25414 15432
rect 25594 15252 25614 15432
rect 25394 15232 25614 15252
rect 25714 15772 26074 15792
rect 25714 15412 25734 15772
rect 26054 15412 26074 15772
rect 26154 15772 26574 17352
rect 26154 15612 26174 15772
rect 26554 15612 26574 15772
rect 26154 15592 26574 15612
rect 26674 17672 26894 17692
rect 26674 17192 26694 17672
rect 26874 17192 26894 17672
rect 25714 15132 26074 15412
rect 26674 15432 26894 17192
rect 27154 16552 27474 17832
rect 27154 16372 27174 16552
rect 27454 16372 27474 16552
rect 27154 16352 27474 16372
rect 27554 18032 27674 18052
rect 27554 17812 27574 18032
rect 27654 17812 27674 18032
rect 27554 16572 27674 17812
rect 27734 17352 27754 18172
rect 27834 17352 27854 18172
rect 27734 17032 27854 17352
rect 27734 16812 27754 17032
rect 27834 16812 27854 17032
rect 27734 16792 27854 16812
rect 27554 16352 27574 16572
rect 27654 16352 27674 16572
rect 26674 15252 26694 15432
rect 26874 15252 26894 15432
rect 27554 16312 27674 16352
rect 27554 15412 27574 16312
rect 27654 15412 27674 16312
rect 27554 15392 27674 15412
rect 26674 15232 26894 15252
rect 25714 14972 25734 15132
rect 26054 14972 26074 15132
rect 25714 14952 26074 14972
rect 24014 14912 24994 14932
rect 2490 2500 2506 2600
rect 2888 2500 2906 2600
rect 2490 2396 2906 2500
rect 29325 1442 29636 19032
rect 26876 1430 29636 1442
rect 26876 1146 26910 1430
rect 27002 1146 29636 1430
rect 26876 1131 29636 1146
<< via3 >>
rect 29480 44480 29580 44600
rect 28740 44280 28860 44400
rect 28000 44040 28120 44200
rect 27240 43820 27400 44000
rect 26520 43620 26660 43760
rect 25760 43420 25940 43540
rect 25020 43220 25200 43340
rect 24280 43000 24460 43140
rect 5676 37418 11236 37938
rect 5676 37198 7436 37418
rect 7436 37198 10666 37418
rect 10666 37198 11236 37418
rect 5676 35848 7446 36078
rect 7446 35848 10656 36078
rect 10656 35848 11256 36078
rect 5676 35258 11256 35848
rect 12976 37158 13356 37978
rect 12536 35218 12856 35578
rect 14556 37158 14636 37978
rect 18464 37536 24024 38056
rect 18464 37316 20224 37536
rect 20224 37316 23454 37536
rect 23454 37316 24024 37536
rect 14376 35218 14456 36118
rect 18464 35966 20234 36196
rect 20234 35966 23444 36196
rect 23444 35966 24044 36196
rect 18464 35376 24044 35966
rect 25764 37276 26144 38096
rect 25324 35336 25644 35696
rect 27344 37276 27424 38096
rect 27164 35336 27244 36236
rect 5696 31492 11256 32012
rect 5696 31272 7456 31492
rect 7456 31272 10686 31492
rect 10686 31272 11256 31492
rect 5696 29922 7466 30152
rect 7466 29922 10676 30152
rect 10676 29922 11276 30152
rect 5696 29332 11276 29922
rect 12996 31232 13376 32052
rect 12556 29292 12876 29652
rect 14576 31232 14656 32052
rect 18428 31416 23988 31936
rect 18428 31196 20188 31416
rect 20188 31196 23418 31416
rect 23418 31196 23988 31416
rect 14396 29292 14476 30192
rect 18428 29846 20198 30076
rect 20198 29846 23408 30076
rect 23408 29846 24008 30076
rect 18428 29256 24008 29846
rect 25728 31156 26108 31976
rect 25288 29216 25608 29576
rect 27308 31156 27388 31976
rect 27128 29216 27208 30116
rect 5816 24788 11376 25308
rect 5816 24568 7576 24788
rect 7576 24568 10806 24788
rect 10806 24568 11376 24788
rect 5816 23218 7586 23448
rect 7586 23218 10796 23448
rect 10796 23218 11396 23448
rect 5816 22628 11396 23218
rect 13116 24528 13496 25348
rect 12676 22588 12996 22948
rect 14696 24528 14776 25348
rect 18524 24658 24084 25178
rect 18524 24438 20284 24658
rect 20284 24438 23514 24658
rect 23514 24438 24084 24658
rect 14516 22588 14596 23488
rect 18524 23088 20294 23318
rect 20294 23088 23504 23318
rect 23504 23088 24104 23318
rect 18524 22498 24104 23088
rect 25824 24398 26204 25218
rect 25384 22458 25704 22818
rect 27404 24398 27484 25218
rect 27224 22458 27304 23358
rect 5692 17742 11252 18262
rect 5692 17522 7452 17742
rect 7452 17522 10682 17742
rect 10682 17522 11252 17742
rect 5692 16172 7462 16402
rect 7462 16172 10672 16402
rect 10672 16172 11272 16402
rect 5692 15582 11272 16172
rect 12992 17482 13372 18302
rect 12552 15542 12872 15902
rect 14572 17482 14652 18302
rect 18874 17612 24434 18132
rect 18874 17392 20634 17612
rect 20634 17392 23864 17612
rect 23864 17392 24434 17612
rect 14392 15542 14472 16442
rect 18874 16042 20644 16272
rect 20644 16042 23854 16272
rect 23854 16042 24454 16272
rect 18874 15452 24454 16042
rect 26174 17352 26554 18172
rect 25734 15412 26054 15772
rect 27754 17352 27834 18172
rect 27574 15412 27654 16312
rect 2506 2500 2888 2600
rect 26910 1146 27002 1430
<< metal4 >>
rect 798 44486 858 45152
rect 1534 44486 1594 45152
rect 2270 44486 2330 45152
rect 3006 44486 3066 45152
rect 3742 44486 3802 45152
rect 4478 44486 4538 45152
rect 5214 44486 5274 45152
rect 5950 44486 6010 45152
rect 6686 44486 6746 45152
rect 7422 44486 7482 45152
rect 8158 44486 8218 45152
rect 8894 44486 8954 45152
rect 9630 44486 9690 45152
rect 10366 44486 10426 45152
rect 11102 44486 11162 45152
rect 11838 44486 11898 45152
rect 12574 44486 12634 45152
rect 13310 44486 13370 45152
rect 14046 44486 14106 45152
rect 14782 44486 14842 45152
rect 15518 44486 15578 45152
rect 16254 44486 16314 45152
rect 16990 44486 17050 45152
rect 17726 44486 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 798 44426 23156 44486
rect 1000 38600 1300 44152
rect 23096 42192 23156 44426
rect 24350 43160 24410 45152
rect 25086 43360 25146 45152
rect 25822 43560 25882 45152
rect 26558 43780 26618 45152
rect 27294 44020 27354 45152
rect 28030 44220 28090 45152
rect 28766 44420 28826 45152
rect 29502 44620 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 29460 44600 29600 44620
rect 29460 44480 29480 44600
rect 29580 44480 29600 44600
rect 29460 44460 29600 44480
rect 28720 44400 28880 44420
rect 28720 44280 28740 44400
rect 28860 44280 28880 44400
rect 28720 44260 28880 44280
rect 27980 44200 28140 44220
rect 27980 44040 28000 44200
rect 28120 44040 28140 44200
rect 27980 44020 28140 44040
rect 27220 44000 27420 44020
rect 27220 43820 27240 44000
rect 27400 43820 27420 44000
rect 27220 43800 27420 43820
rect 26500 43760 26680 43780
rect 26500 43620 26520 43760
rect 26660 43620 26680 43760
rect 26500 43600 26680 43620
rect 25720 43540 25960 43560
rect 25720 43420 25760 43540
rect 25940 43420 25960 43540
rect 25720 43400 25960 43420
rect 25000 43340 25220 43360
rect 25000 43220 25020 43340
rect 25200 43220 25220 43340
rect 25000 43200 25220 43220
rect 24260 43140 24480 43160
rect 24260 43000 24280 43140
rect 24460 43000 24480 43140
rect 24260 42980 24480 43000
rect 31506 42192 31806 44152
rect 23096 42132 31806 42192
rect 1000 38096 28800 38600
rect 1000 38056 25764 38096
rect 1000 37978 18464 38056
rect 1000 37938 12976 37978
rect 1000 37198 5676 37938
rect 11236 37198 12976 37938
rect 1000 37158 12976 37198
rect 13356 37158 14556 37978
rect 14636 37316 18464 37978
rect 24024 37316 25764 38056
rect 14636 37276 25764 37316
rect 26144 37276 27344 38096
rect 27424 37276 28800 38096
rect 14636 37158 28800 37276
rect 1000 37000 28800 37158
rect 1000 32600 1300 37000
rect 31506 36400 31806 42132
rect 5400 36236 31806 36400
rect 5400 36196 27164 36236
rect 5400 36118 18464 36196
rect 5400 36078 14376 36118
rect 5400 35258 5676 36078
rect 11256 35578 14376 36078
rect 11256 35258 12536 35578
rect 5400 35218 12536 35258
rect 12856 35218 14376 35578
rect 14456 35376 18464 36118
rect 24044 35696 27164 36196
rect 24044 35376 25324 35696
rect 14456 35336 25324 35376
rect 25644 35336 27164 35696
rect 27244 35336 31806 36236
rect 14456 35218 31806 35336
rect 5400 35000 31806 35218
rect 1000 32052 28800 32600
rect 1000 32012 12996 32052
rect 1000 31272 5696 32012
rect 11256 31272 12996 32012
rect 1000 31232 12996 31272
rect 13376 31232 14576 32052
rect 14656 31976 28800 32052
rect 14656 31936 25728 31976
rect 14656 31232 18428 31936
rect 1000 31196 18428 31232
rect 23988 31196 25728 31936
rect 1000 31156 25728 31196
rect 26108 31156 27308 31976
rect 27388 31156 28800 31976
rect 1000 31000 28800 31156
rect 1000 25600 1300 31000
rect 31506 30400 31806 35000
rect 5400 30192 31806 30400
rect 5400 30152 14396 30192
rect 5400 29332 5696 30152
rect 11276 29652 14396 30152
rect 11276 29332 12556 29652
rect 5400 29292 12556 29332
rect 12876 29292 14396 29652
rect 14476 30116 31806 30192
rect 14476 30076 27128 30116
rect 14476 29292 18428 30076
rect 5400 29256 18428 29292
rect 24008 29576 27128 30076
rect 24008 29256 25288 29576
rect 5400 29216 25288 29256
rect 25608 29216 27128 29576
rect 27208 29216 31806 30116
rect 5400 29000 31806 29216
rect 1000 25348 28800 25600
rect 1000 25308 13116 25348
rect 1000 24568 5816 25308
rect 11376 24568 13116 25308
rect 1000 24528 13116 24568
rect 13496 24528 14696 25348
rect 14776 25218 28800 25348
rect 14776 25178 25824 25218
rect 14776 24528 18524 25178
rect 1000 24438 18524 24528
rect 24084 24438 25824 25178
rect 1000 24398 25824 24438
rect 26204 24398 27404 25218
rect 27484 24398 28800 25218
rect 1000 24000 28800 24398
rect 1000 18400 1300 24000
rect 31506 23600 31806 29000
rect 5400 23488 31806 23600
rect 5400 23448 14516 23488
rect 5400 22628 5816 23448
rect 11396 22948 14516 23448
rect 11396 22628 12676 22948
rect 5400 22588 12676 22628
rect 12996 22588 14516 22948
rect 14596 23358 31806 23488
rect 14596 23318 27224 23358
rect 14596 22588 18524 23318
rect 5400 22498 18524 22588
rect 24104 22818 27224 23318
rect 24104 22498 25384 22818
rect 5400 22458 25384 22498
rect 25704 22458 27224 22818
rect 27304 22458 31806 23358
rect 5400 22200 31806 22458
rect 1000 18302 28800 18400
rect 1000 18262 12992 18302
rect 1000 17522 5692 18262
rect 11252 17522 12992 18262
rect 1000 17482 12992 17522
rect 13372 17482 14572 18302
rect 14652 18172 28800 18302
rect 14652 18132 26174 18172
rect 14652 17482 18874 18132
rect 1000 17392 18874 17482
rect 24434 17392 26174 18132
rect 1000 17352 26174 17392
rect 26554 17352 27754 18172
rect 27834 17352 28800 18172
rect 1000 17200 28800 17352
rect 1000 1000 1300 17200
rect 31506 16800 31806 22200
rect 5400 16442 31806 16800
rect 5400 16402 14392 16442
rect 5400 15582 5692 16402
rect 11272 15902 14392 16402
rect 11272 15582 12552 15902
rect 5400 15542 12552 15582
rect 12872 15542 14392 15902
rect 14472 16312 31806 16442
rect 14472 16272 27574 16312
rect 14472 15542 18874 16272
rect 5400 15452 18874 15542
rect 24454 15772 27574 16272
rect 24454 15452 25734 15772
rect 5400 15412 25734 15452
rect 26054 15412 27574 15772
rect 27654 15412 31806 16312
rect 5400 15400 31806 15412
rect 18814 15392 28394 15400
rect 2417 2600 28525 2609
rect 2417 2500 2506 2600
rect 2888 2500 28525 2600
rect 2417 2491 28525 2500
rect 26896 1430 27016 1456
rect 26896 1146 26910 1430
rect 27002 1146 27016 1430
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 200
rect 13648 0 13768 200
rect 18064 0 18184 200
rect 22480 0 22600 200
rect 26896 0 27016 1146
rect 28407 482 28525 2491
rect 31506 1000 31806 15400
rect 28406 362 31432 482
rect 31312 0 31432 362
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 31506 1000 31806 44152 1 FreeSans 200 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 1000 1000 1300 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal3 25714 18832 26074 19352 0 FreeSans 1600 0 0 0 distortionUnit_7.CTRL
flabel via3 18874 15452 24454 16272 0 FreeSans 1600 0 0 0 distortionUnit_7.VSS
flabel via3 18874 17392 24434 18132 0 FreeSans 1600 0 0 0 distortionUnit_7.VDD
flabel metal3 27154 18012 27474 19352 0 FreeSans 1600 0 0 0 distortionUnit_7.OUT
flabel metal3 18354 18492 18694 19212 0 FreeSans 1600 0 0 0 distortionUnit_7.IN
flabel metal2 25594 16832 25914 17052 0 FreeSans 1600 0 0 0 distortionUnit_7.tgate_1.IN
flabel metal2 25594 16352 25914 16572 0 FreeSans 1600 0 0 0 distortionUnit_7.tgate_1.OUT
flabel metal2 25594 17172 26134 17392 0 FreeSans 1600 0 0 0 distortionUnit_7.tgate_1.CTRLB
flabel metal2 25594 16012 26134 16232 0 FreeSans 1600 0 0 0 distortionUnit_7.tgate_1.CTRL
flabel metal1 26954 16832 27274 17052 0 FreeSans 1600 0 0 0 distortionUnit_7.tgate_1.VDD
flabel metal1 26954 16352 27274 16572 0 FreeSans 1600 0 0 0 distortionUnit_7.tgate_1.VSS
flabel metal2 25594 18292 25914 18512 0 FreeSans 1600 0 0 0 distortionUnit_7.tgate_0.IN
flabel metal2 25594 17812 25914 18032 0 FreeSans 1600 0 0 0 distortionUnit_7.tgate_0.OUT
flabel metal2 25594 18632 26134 18852 0 FreeSans 1600 0 0 0 distortionUnit_7.tgate_0.CTRLB
flabel metal2 25594 17472 26134 17692 0 FreeSans 1600 0 0 0 distortionUnit_7.tgate_0.CTRL
flabel metal1 26954 18292 27274 18512 0 FreeSans 1600 0 0 0 distortionUnit_7.tgate_0.VDD
flabel metal1 26954 17812 27274 18032 0 FreeSans 1600 0 0 0 distortionUnit_7.tgate_0.VSS
flabel metal1 26599 15086 26647 15112 0 FreeSans 200 0 0 0 distortionUnit_7.sky130_fd_sc_hd__tap_2_0.VGND
flabel metal1 26601 15633 26655 15655 0 FreeSans 200 0 0 0 distortionUnit_7.sky130_fd_sc_hd__tap_2_0.VPWR
flabel locali 26615 15531 26640 15556 0 FreeSans 250 0 0 0 distortionUnit_7.sky130_fd_sc_hd__tap_2_0.VPB
flabel locali 26700 15192 26735 15222 0 FreeSans 250 0 0 0 distortionUnit_7.sky130_fd_sc_hd__tap_2_0.VNB
flabel locali 26708 15525 26730 15554 0 FreeSans 250 0 0 0 distortionUnit_7.sky130_fd_sc_hd__tap_2_0.VPB
rlabel comment 26580 15100 26580 15100 4 distortionUnit_7.sky130_fd_sc_hd__tap_2_0.tap_2
rlabel metal1 26580 15052 26764 15148 1 distortionUnit_7.sky130_fd_sc_hd__tap_2_0.VGND
rlabel metal1 26580 15596 26764 15692 1 distortionUnit_7.sky130_fd_sc_hd__tap_2_0.VPWR
flabel locali 25965 15321 25999 15355 0 FreeSans 250 0 0 0 distortionUnit_7.sky130_fd_sc_hd__inv_8_0.A
flabel locali 26057 15321 26091 15355 0 FreeSans 250 0 0 0 distortionUnit_7.sky130_fd_sc_hd__inv_8_0.A
flabel locali 26149 15321 26183 15355 0 FreeSans 250 0 0 0 distortionUnit_7.sky130_fd_sc_hd__inv_8_0.A
flabel locali 26241 15321 26275 15355 0 FreeSans 250 0 0 0 distortionUnit_7.sky130_fd_sc_hd__inv_8_0.A
flabel locali 26333 15321 26367 15355 0 FreeSans 250 0 0 0 distortionUnit_7.sky130_fd_sc_hd__inv_8_0.A
flabel locali 26425 15321 26459 15355 0 FreeSans 250 0 0 0 distortionUnit_7.sky130_fd_sc_hd__inv_8_0.A
flabel locali 26517 15321 26551 15355 0 FreeSans 250 0 0 0 distortionUnit_7.sky130_fd_sc_hd__inv_8_0.Y
flabel locali 25781 15321 25815 15355 0 FreeSans 250 0 0 0 distortionUnit_7.sky130_fd_sc_hd__inv_8_0.Y
flabel pwell 25781 15083 25815 15117 0 FreeSans 200 0 0 0 distortionUnit_7.sky130_fd_sc_hd__inv_8_0.VNB
flabel nwell 25781 15627 25815 15661 0 FreeSans 200 0 0 0 distortionUnit_7.sky130_fd_sc_hd__inv_8_0.VPB
flabel metal1 25781 15083 25815 15117 0 FreeSans 200 0 0 0 distortionUnit_7.sky130_fd_sc_hd__inv_8_0.VGND
flabel metal1 25781 15627 25815 15661 0 FreeSans 200 0 0 0 distortionUnit_7.sky130_fd_sc_hd__inv_8_0.VPWR
rlabel comment 25752 15100 25752 15100 4 distortionUnit_7.sky130_fd_sc_hd__inv_8_0.inv_8
rlabel metal1 25752 15052 26580 15148 1 distortionUnit_7.sky130_fd_sc_hd__inv_8_0.VGND
rlabel metal1 25752 15596 26580 15692 1 distortionUnit_7.sky130_fd_sc_hd__inv_8_0.VPWR
flabel metal3 23434 16652 23824 17042 0 FreeSans 800 0 0 0 distortionUnit_7.myOpamp_0.INn
flabel metal3 21404 16942 23064 17192 0 FreeSans 800 0 0 0 distortionUnit_7.myOpamp_0.OUT
flabel metal3 20644 16042 23854 16292 0 FreeSans 800 0 0 0 distortionUnit_7.myOpamp_0.VSS
flabel metal3 20634 17342 23864 17612 0 FreeSans 800 0 0 0 distortionUnit_7.myOpamp_0.VDD
flabel metal3 20674 16942 21064 17252 0 FreeSans 800 0 0 0 distortionUnit_7.myOpamp_0.INp
flabel metal3 25364 25878 25724 26398 0 FreeSans 1600 0 0 0 distortionUnit_6.CTRL
flabel via3 18524 22498 24104 23318 0 FreeSans 1600 0 0 0 distortionUnit_6.VSS
flabel via3 18524 24438 24084 25178 0 FreeSans 1600 0 0 0 distortionUnit_6.VDD
flabel metal3 26804 25058 27124 26398 0 FreeSans 1600 0 0 0 distortionUnit_6.OUT
flabel metal3 18004 25538 18344 26258 0 FreeSans 1600 0 0 0 distortionUnit_6.IN
flabel metal2 25244 23878 25564 24098 0 FreeSans 1600 0 0 0 distortionUnit_6.tgate_1.IN
flabel metal2 25244 23398 25564 23618 0 FreeSans 1600 0 0 0 distortionUnit_6.tgate_1.OUT
flabel metal2 25244 24218 25784 24438 0 FreeSans 1600 0 0 0 distortionUnit_6.tgate_1.CTRLB
flabel metal2 25244 23058 25784 23278 0 FreeSans 1600 0 0 0 distortionUnit_6.tgate_1.CTRL
flabel metal1 26604 23878 26924 24098 0 FreeSans 1600 0 0 0 distortionUnit_6.tgate_1.VDD
flabel metal1 26604 23398 26924 23618 0 FreeSans 1600 0 0 0 distortionUnit_6.tgate_1.VSS
flabel metal2 25244 25338 25564 25558 0 FreeSans 1600 0 0 0 distortionUnit_6.tgate_0.IN
flabel metal2 25244 24858 25564 25078 0 FreeSans 1600 0 0 0 distortionUnit_6.tgate_0.OUT
flabel metal2 25244 25678 25784 25898 0 FreeSans 1600 0 0 0 distortionUnit_6.tgate_0.CTRLB
flabel metal2 25244 24518 25784 24738 0 FreeSans 1600 0 0 0 distortionUnit_6.tgate_0.CTRL
flabel metal1 26604 25338 26924 25558 0 FreeSans 1600 0 0 0 distortionUnit_6.tgate_0.VDD
flabel metal1 26604 24858 26924 25078 0 FreeSans 1600 0 0 0 distortionUnit_6.tgate_0.VSS
flabel metal1 26249 22132 26297 22158 0 FreeSans 200 0 0 0 distortionUnit_6.sky130_fd_sc_hd__tap_2_0.VGND
flabel metal1 26251 22679 26305 22701 0 FreeSans 200 0 0 0 distortionUnit_6.sky130_fd_sc_hd__tap_2_0.VPWR
flabel locali 26265 22577 26290 22602 0 FreeSans 250 0 0 0 distortionUnit_6.sky130_fd_sc_hd__tap_2_0.VPB
flabel locali 26350 22238 26385 22268 0 FreeSans 250 0 0 0 distortionUnit_6.sky130_fd_sc_hd__tap_2_0.VNB
flabel locali 26358 22571 26380 22600 0 FreeSans 250 0 0 0 distortionUnit_6.sky130_fd_sc_hd__tap_2_0.VPB
rlabel comment 26230 22146 26230 22146 4 distortionUnit_6.sky130_fd_sc_hd__tap_2_0.tap_2
rlabel metal1 26230 22098 26414 22194 1 distortionUnit_6.sky130_fd_sc_hd__tap_2_0.VGND
rlabel metal1 26230 22642 26414 22738 1 distortionUnit_6.sky130_fd_sc_hd__tap_2_0.VPWR
flabel locali 25615 22367 25649 22401 0 FreeSans 250 0 0 0 distortionUnit_6.sky130_fd_sc_hd__inv_8_0.A
flabel locali 25707 22367 25741 22401 0 FreeSans 250 0 0 0 distortionUnit_6.sky130_fd_sc_hd__inv_8_0.A
flabel locali 25799 22367 25833 22401 0 FreeSans 250 0 0 0 distortionUnit_6.sky130_fd_sc_hd__inv_8_0.A
flabel locali 25891 22367 25925 22401 0 FreeSans 250 0 0 0 distortionUnit_6.sky130_fd_sc_hd__inv_8_0.A
flabel locali 25983 22367 26017 22401 0 FreeSans 250 0 0 0 distortionUnit_6.sky130_fd_sc_hd__inv_8_0.A
flabel locali 26075 22367 26109 22401 0 FreeSans 250 0 0 0 distortionUnit_6.sky130_fd_sc_hd__inv_8_0.A
flabel locali 26167 22367 26201 22401 0 FreeSans 250 0 0 0 distortionUnit_6.sky130_fd_sc_hd__inv_8_0.Y
flabel locali 25431 22367 25465 22401 0 FreeSans 250 0 0 0 distortionUnit_6.sky130_fd_sc_hd__inv_8_0.Y
flabel pwell 25431 22129 25465 22163 0 FreeSans 200 0 0 0 distortionUnit_6.sky130_fd_sc_hd__inv_8_0.VNB
flabel nwell 25431 22673 25465 22707 0 FreeSans 200 0 0 0 distortionUnit_6.sky130_fd_sc_hd__inv_8_0.VPB
flabel metal1 25431 22129 25465 22163 0 FreeSans 200 0 0 0 distortionUnit_6.sky130_fd_sc_hd__inv_8_0.VGND
flabel metal1 25431 22673 25465 22707 0 FreeSans 200 0 0 0 distortionUnit_6.sky130_fd_sc_hd__inv_8_0.VPWR
rlabel comment 25402 22146 25402 22146 4 distortionUnit_6.sky130_fd_sc_hd__inv_8_0.inv_8
rlabel metal1 25402 22098 26230 22194 1 distortionUnit_6.sky130_fd_sc_hd__inv_8_0.VGND
rlabel metal1 25402 22642 26230 22738 1 distortionUnit_6.sky130_fd_sc_hd__inv_8_0.VPWR
flabel metal3 23084 23698 23474 24088 0 FreeSans 800 0 0 0 distortionUnit_6.myOpamp_0.INn
flabel metal3 21054 23988 22714 24238 0 FreeSans 800 0 0 0 distortionUnit_6.myOpamp_0.OUT
flabel metal3 20294 23088 23504 23338 0 FreeSans 800 0 0 0 distortionUnit_6.myOpamp_0.VSS
flabel metal3 20284 24388 23514 24658 0 FreeSans 800 0 0 0 distortionUnit_6.myOpamp_0.VDD
flabel metal3 20324 23988 20714 24298 0 FreeSans 800 0 0 0 distortionUnit_6.myOpamp_0.INp
flabel metal3 12656 26008 13016 26528 0 FreeSans 1600 0 0 0 distortionUnit_5.CTRL
flabel via3 5816 22628 11396 23448 0 FreeSans 1600 0 0 0 distortionUnit_5.VSS
flabel via3 5816 24568 11376 25308 0 FreeSans 1600 0 0 0 distortionUnit_5.VDD
flabel metal3 14096 25188 14416 26528 0 FreeSans 1600 0 0 0 distortionUnit_5.OUT
flabel metal3 5296 25668 5636 26388 0 FreeSans 1600 0 0 0 distortionUnit_5.IN
flabel metal2 12536 24008 12856 24228 0 FreeSans 1600 0 0 0 distortionUnit_5.tgate_1.IN
flabel metal2 12536 23528 12856 23748 0 FreeSans 1600 0 0 0 distortionUnit_5.tgate_1.OUT
flabel metal2 12536 24348 13076 24568 0 FreeSans 1600 0 0 0 distortionUnit_5.tgate_1.CTRLB
flabel metal2 12536 23188 13076 23408 0 FreeSans 1600 0 0 0 distortionUnit_5.tgate_1.CTRL
flabel metal1 13896 24008 14216 24228 0 FreeSans 1600 0 0 0 distortionUnit_5.tgate_1.VDD
flabel metal1 13896 23528 14216 23748 0 FreeSans 1600 0 0 0 distortionUnit_5.tgate_1.VSS
flabel metal2 12536 25468 12856 25688 0 FreeSans 1600 0 0 0 distortionUnit_5.tgate_0.IN
flabel metal2 12536 24988 12856 25208 0 FreeSans 1600 0 0 0 distortionUnit_5.tgate_0.OUT
flabel metal2 12536 25808 13076 26028 0 FreeSans 1600 0 0 0 distortionUnit_5.tgate_0.CTRLB
flabel metal2 12536 24648 13076 24868 0 FreeSans 1600 0 0 0 distortionUnit_5.tgate_0.CTRL
flabel metal1 13896 25468 14216 25688 0 FreeSans 1600 0 0 0 distortionUnit_5.tgate_0.VDD
flabel metal1 13896 24988 14216 25208 0 FreeSans 1600 0 0 0 distortionUnit_5.tgate_0.VSS
flabel metal1 13541 22262 13589 22288 0 FreeSans 200 0 0 0 distortionUnit_5.sky130_fd_sc_hd__tap_2_0.VGND
flabel metal1 13543 22809 13597 22831 0 FreeSans 200 0 0 0 distortionUnit_5.sky130_fd_sc_hd__tap_2_0.VPWR
flabel locali 13557 22707 13582 22732 0 FreeSans 250 0 0 0 distortionUnit_5.sky130_fd_sc_hd__tap_2_0.VPB
flabel locali 13642 22368 13677 22398 0 FreeSans 250 0 0 0 distortionUnit_5.sky130_fd_sc_hd__tap_2_0.VNB
flabel locali 13650 22701 13672 22730 0 FreeSans 250 0 0 0 distortionUnit_5.sky130_fd_sc_hd__tap_2_0.VPB
rlabel comment 13522 22276 13522 22276 4 distortionUnit_5.sky130_fd_sc_hd__tap_2_0.tap_2
rlabel metal1 13522 22228 13706 22324 1 distortionUnit_5.sky130_fd_sc_hd__tap_2_0.VGND
rlabel metal1 13522 22772 13706 22868 1 distortionUnit_5.sky130_fd_sc_hd__tap_2_0.VPWR
flabel locali 12907 22497 12941 22531 0 FreeSans 250 0 0 0 distortionUnit_5.sky130_fd_sc_hd__inv_8_0.A
flabel locali 12999 22497 13033 22531 0 FreeSans 250 0 0 0 distortionUnit_5.sky130_fd_sc_hd__inv_8_0.A
flabel locali 13091 22497 13125 22531 0 FreeSans 250 0 0 0 distortionUnit_5.sky130_fd_sc_hd__inv_8_0.A
flabel locali 13183 22497 13217 22531 0 FreeSans 250 0 0 0 distortionUnit_5.sky130_fd_sc_hd__inv_8_0.A
flabel locali 13275 22497 13309 22531 0 FreeSans 250 0 0 0 distortionUnit_5.sky130_fd_sc_hd__inv_8_0.A
flabel locali 13367 22497 13401 22531 0 FreeSans 250 0 0 0 distortionUnit_5.sky130_fd_sc_hd__inv_8_0.A
flabel locali 13459 22497 13493 22531 0 FreeSans 250 0 0 0 distortionUnit_5.sky130_fd_sc_hd__inv_8_0.Y
flabel locali 12723 22497 12757 22531 0 FreeSans 250 0 0 0 distortionUnit_5.sky130_fd_sc_hd__inv_8_0.Y
flabel pwell 12723 22259 12757 22293 0 FreeSans 200 0 0 0 distortionUnit_5.sky130_fd_sc_hd__inv_8_0.VNB
flabel nwell 12723 22803 12757 22837 0 FreeSans 200 0 0 0 distortionUnit_5.sky130_fd_sc_hd__inv_8_0.VPB
flabel metal1 12723 22259 12757 22293 0 FreeSans 200 0 0 0 distortionUnit_5.sky130_fd_sc_hd__inv_8_0.VGND
flabel metal1 12723 22803 12757 22837 0 FreeSans 200 0 0 0 distortionUnit_5.sky130_fd_sc_hd__inv_8_0.VPWR
rlabel comment 12694 22276 12694 22276 4 distortionUnit_5.sky130_fd_sc_hd__inv_8_0.inv_8
rlabel metal1 12694 22228 13522 22324 1 distortionUnit_5.sky130_fd_sc_hd__inv_8_0.VGND
rlabel metal1 12694 22772 13522 22868 1 distortionUnit_5.sky130_fd_sc_hd__inv_8_0.VPWR
flabel metal3 10376 23828 10766 24218 0 FreeSans 800 0 0 0 distortionUnit_5.myOpamp_0.INn
flabel metal3 8346 24118 10006 24368 0 FreeSans 800 0 0 0 distortionUnit_5.myOpamp_0.OUT
flabel metal3 7586 23218 10796 23468 0 FreeSans 800 0 0 0 distortionUnit_5.myOpamp_0.VSS
flabel metal3 7576 24518 10806 24788 0 FreeSans 800 0 0 0 distortionUnit_5.myOpamp_0.VDD
flabel metal3 7616 24118 8006 24428 0 FreeSans 800 0 0 0 distortionUnit_5.myOpamp_0.INp
flabel metal3 25268 32636 25628 33156 0 FreeSans 1600 0 0 0 distortionUnit_4.CTRL
flabel via3 18428 29256 24008 30076 0 FreeSans 1600 0 0 0 distortionUnit_4.VSS
flabel via3 18428 31196 23988 31936 0 FreeSans 1600 0 0 0 distortionUnit_4.VDD
flabel metal3 26708 31816 27028 33156 0 FreeSans 1600 0 0 0 distortionUnit_4.OUT
flabel metal3 17908 32296 18248 33016 0 FreeSans 1600 0 0 0 distortionUnit_4.IN
flabel metal2 25148 30636 25468 30856 0 FreeSans 1600 0 0 0 distortionUnit_4.tgate_1.IN
flabel metal2 25148 30156 25468 30376 0 FreeSans 1600 0 0 0 distortionUnit_4.tgate_1.OUT
flabel metal2 25148 30976 25688 31196 0 FreeSans 1600 0 0 0 distortionUnit_4.tgate_1.CTRLB
flabel metal2 25148 29816 25688 30036 0 FreeSans 1600 0 0 0 distortionUnit_4.tgate_1.CTRL
flabel metal1 26508 30636 26828 30856 0 FreeSans 1600 0 0 0 distortionUnit_4.tgate_1.VDD
flabel metal1 26508 30156 26828 30376 0 FreeSans 1600 0 0 0 distortionUnit_4.tgate_1.VSS
flabel metal2 25148 32096 25468 32316 0 FreeSans 1600 0 0 0 distortionUnit_4.tgate_0.IN
flabel metal2 25148 31616 25468 31836 0 FreeSans 1600 0 0 0 distortionUnit_4.tgate_0.OUT
flabel metal2 25148 32436 25688 32656 0 FreeSans 1600 0 0 0 distortionUnit_4.tgate_0.CTRLB
flabel metal2 25148 31276 25688 31496 0 FreeSans 1600 0 0 0 distortionUnit_4.tgate_0.CTRL
flabel metal1 26508 32096 26828 32316 0 FreeSans 1600 0 0 0 distortionUnit_4.tgate_0.VDD
flabel metal1 26508 31616 26828 31836 0 FreeSans 1600 0 0 0 distortionUnit_4.tgate_0.VSS
flabel metal1 26153 28890 26201 28916 0 FreeSans 200 0 0 0 distortionUnit_4.sky130_fd_sc_hd__tap_2_0.VGND
flabel metal1 26155 29437 26209 29459 0 FreeSans 200 0 0 0 distortionUnit_4.sky130_fd_sc_hd__tap_2_0.VPWR
flabel locali 26169 29335 26194 29360 0 FreeSans 250 0 0 0 distortionUnit_4.sky130_fd_sc_hd__tap_2_0.VPB
flabel locali 26254 28996 26289 29026 0 FreeSans 250 0 0 0 distortionUnit_4.sky130_fd_sc_hd__tap_2_0.VNB
flabel locali 26262 29329 26284 29358 0 FreeSans 250 0 0 0 distortionUnit_4.sky130_fd_sc_hd__tap_2_0.VPB
rlabel comment 26134 28904 26134 28904 4 distortionUnit_4.sky130_fd_sc_hd__tap_2_0.tap_2
rlabel metal1 26134 28856 26318 28952 1 distortionUnit_4.sky130_fd_sc_hd__tap_2_0.VGND
rlabel metal1 26134 29400 26318 29496 1 distortionUnit_4.sky130_fd_sc_hd__tap_2_0.VPWR
flabel locali 25519 29125 25553 29159 0 FreeSans 250 0 0 0 distortionUnit_4.sky130_fd_sc_hd__inv_8_0.A
flabel locali 25611 29125 25645 29159 0 FreeSans 250 0 0 0 distortionUnit_4.sky130_fd_sc_hd__inv_8_0.A
flabel locali 25703 29125 25737 29159 0 FreeSans 250 0 0 0 distortionUnit_4.sky130_fd_sc_hd__inv_8_0.A
flabel locali 25795 29125 25829 29159 0 FreeSans 250 0 0 0 distortionUnit_4.sky130_fd_sc_hd__inv_8_0.A
flabel locali 25887 29125 25921 29159 0 FreeSans 250 0 0 0 distortionUnit_4.sky130_fd_sc_hd__inv_8_0.A
flabel locali 25979 29125 26013 29159 0 FreeSans 250 0 0 0 distortionUnit_4.sky130_fd_sc_hd__inv_8_0.A
flabel locali 26071 29125 26105 29159 0 FreeSans 250 0 0 0 distortionUnit_4.sky130_fd_sc_hd__inv_8_0.Y
flabel locali 25335 29125 25369 29159 0 FreeSans 250 0 0 0 distortionUnit_4.sky130_fd_sc_hd__inv_8_0.Y
flabel pwell 25335 28887 25369 28921 0 FreeSans 200 0 0 0 distortionUnit_4.sky130_fd_sc_hd__inv_8_0.VNB
flabel nwell 25335 29431 25369 29465 0 FreeSans 200 0 0 0 distortionUnit_4.sky130_fd_sc_hd__inv_8_0.VPB
flabel metal1 25335 28887 25369 28921 0 FreeSans 200 0 0 0 distortionUnit_4.sky130_fd_sc_hd__inv_8_0.VGND
flabel metal1 25335 29431 25369 29465 0 FreeSans 200 0 0 0 distortionUnit_4.sky130_fd_sc_hd__inv_8_0.VPWR
rlabel comment 25306 28904 25306 28904 4 distortionUnit_4.sky130_fd_sc_hd__inv_8_0.inv_8
rlabel metal1 25306 28856 26134 28952 1 distortionUnit_4.sky130_fd_sc_hd__inv_8_0.VGND
rlabel metal1 25306 29400 26134 29496 1 distortionUnit_4.sky130_fd_sc_hd__inv_8_0.VPWR
flabel metal3 22988 30456 23378 30846 0 FreeSans 800 0 0 0 distortionUnit_4.myOpamp_0.INn
flabel metal3 20958 30746 22618 30996 0 FreeSans 800 0 0 0 distortionUnit_4.myOpamp_0.OUT
flabel metal3 20198 29846 23408 30096 0 FreeSans 800 0 0 0 distortionUnit_4.myOpamp_0.VSS
flabel metal3 20188 31146 23418 31416 0 FreeSans 800 0 0 0 distortionUnit_4.myOpamp_0.VDD
flabel metal3 20228 30746 20618 31056 0 FreeSans 800 0 0 0 distortionUnit_4.myOpamp_0.INp
flabel metal3 12536 32712 12896 33232 0 FreeSans 1600 0 0 0 distortionUnit_3.CTRL
flabel via3 5696 29332 11276 30152 0 FreeSans 1600 0 0 0 distortionUnit_3.VSS
flabel via3 5696 31272 11256 32012 0 FreeSans 1600 0 0 0 distortionUnit_3.VDD
flabel metal3 13976 31892 14296 33232 0 FreeSans 1600 0 0 0 distortionUnit_3.OUT
flabel metal3 5176 32372 5516 33092 0 FreeSans 1600 0 0 0 distortionUnit_3.IN
flabel metal2 12416 30712 12736 30932 0 FreeSans 1600 0 0 0 distortionUnit_3.tgate_1.IN
flabel metal2 12416 30232 12736 30452 0 FreeSans 1600 0 0 0 distortionUnit_3.tgate_1.OUT
flabel metal2 12416 31052 12956 31272 0 FreeSans 1600 0 0 0 distortionUnit_3.tgate_1.CTRLB
flabel metal2 12416 29892 12956 30112 0 FreeSans 1600 0 0 0 distortionUnit_3.tgate_1.CTRL
flabel metal1 13776 30712 14096 30932 0 FreeSans 1600 0 0 0 distortionUnit_3.tgate_1.VDD
flabel metal1 13776 30232 14096 30452 0 FreeSans 1600 0 0 0 distortionUnit_3.tgate_1.VSS
flabel metal2 12416 32172 12736 32392 0 FreeSans 1600 0 0 0 distortionUnit_3.tgate_0.IN
flabel metal2 12416 31692 12736 31912 0 FreeSans 1600 0 0 0 distortionUnit_3.tgate_0.OUT
flabel metal2 12416 32512 12956 32732 0 FreeSans 1600 0 0 0 distortionUnit_3.tgate_0.CTRLB
flabel metal2 12416 31352 12956 31572 0 FreeSans 1600 0 0 0 distortionUnit_3.tgate_0.CTRL
flabel metal1 13776 32172 14096 32392 0 FreeSans 1600 0 0 0 distortionUnit_3.tgate_0.VDD
flabel metal1 13776 31692 14096 31912 0 FreeSans 1600 0 0 0 distortionUnit_3.tgate_0.VSS
flabel metal1 13421 28966 13469 28992 0 FreeSans 200 0 0 0 distortionUnit_3.sky130_fd_sc_hd__tap_2_0.VGND
flabel metal1 13423 29513 13477 29535 0 FreeSans 200 0 0 0 distortionUnit_3.sky130_fd_sc_hd__tap_2_0.VPWR
flabel locali 13437 29411 13462 29436 0 FreeSans 250 0 0 0 distortionUnit_3.sky130_fd_sc_hd__tap_2_0.VPB
flabel locali 13522 29072 13557 29102 0 FreeSans 250 0 0 0 distortionUnit_3.sky130_fd_sc_hd__tap_2_0.VNB
flabel locali 13530 29405 13552 29434 0 FreeSans 250 0 0 0 distortionUnit_3.sky130_fd_sc_hd__tap_2_0.VPB
rlabel comment 13402 28980 13402 28980 4 distortionUnit_3.sky130_fd_sc_hd__tap_2_0.tap_2
rlabel metal1 13402 28932 13586 29028 1 distortionUnit_3.sky130_fd_sc_hd__tap_2_0.VGND
rlabel metal1 13402 29476 13586 29572 1 distortionUnit_3.sky130_fd_sc_hd__tap_2_0.VPWR
flabel locali 12787 29201 12821 29235 0 FreeSans 250 0 0 0 distortionUnit_3.sky130_fd_sc_hd__inv_8_0.A
flabel locali 12879 29201 12913 29235 0 FreeSans 250 0 0 0 distortionUnit_3.sky130_fd_sc_hd__inv_8_0.A
flabel locali 12971 29201 13005 29235 0 FreeSans 250 0 0 0 distortionUnit_3.sky130_fd_sc_hd__inv_8_0.A
flabel locali 13063 29201 13097 29235 0 FreeSans 250 0 0 0 distortionUnit_3.sky130_fd_sc_hd__inv_8_0.A
flabel locali 13155 29201 13189 29235 0 FreeSans 250 0 0 0 distortionUnit_3.sky130_fd_sc_hd__inv_8_0.A
flabel locali 13247 29201 13281 29235 0 FreeSans 250 0 0 0 distortionUnit_3.sky130_fd_sc_hd__inv_8_0.A
flabel locali 13339 29201 13373 29235 0 FreeSans 250 0 0 0 distortionUnit_3.sky130_fd_sc_hd__inv_8_0.Y
flabel locali 12603 29201 12637 29235 0 FreeSans 250 0 0 0 distortionUnit_3.sky130_fd_sc_hd__inv_8_0.Y
flabel pwell 12603 28963 12637 28997 0 FreeSans 200 0 0 0 distortionUnit_3.sky130_fd_sc_hd__inv_8_0.VNB
flabel nwell 12603 29507 12637 29541 0 FreeSans 200 0 0 0 distortionUnit_3.sky130_fd_sc_hd__inv_8_0.VPB
flabel metal1 12603 28963 12637 28997 0 FreeSans 200 0 0 0 distortionUnit_3.sky130_fd_sc_hd__inv_8_0.VGND
flabel metal1 12603 29507 12637 29541 0 FreeSans 200 0 0 0 distortionUnit_3.sky130_fd_sc_hd__inv_8_0.VPWR
rlabel comment 12574 28980 12574 28980 4 distortionUnit_3.sky130_fd_sc_hd__inv_8_0.inv_8
rlabel metal1 12574 28932 13402 29028 1 distortionUnit_3.sky130_fd_sc_hd__inv_8_0.VGND
rlabel metal1 12574 29476 13402 29572 1 distortionUnit_3.sky130_fd_sc_hd__inv_8_0.VPWR
flabel metal3 10256 30532 10646 30922 0 FreeSans 800 0 0 0 distortionUnit_3.myOpamp_0.INn
flabel metal3 8226 30822 9886 31072 0 FreeSans 800 0 0 0 distortionUnit_3.myOpamp_0.OUT
flabel metal3 7466 29922 10676 30172 0 FreeSans 800 0 0 0 distortionUnit_3.myOpamp_0.VSS
flabel metal3 7456 31222 10686 31492 0 FreeSans 800 0 0 0 distortionUnit_3.myOpamp_0.VDD
flabel metal3 7496 30822 7886 31132 0 FreeSans 800 0 0 0 distortionUnit_3.myOpamp_0.INp
flabel metal3 25304 38756 25664 39276 0 FreeSans 1600 0 0 0 distortionUnit_2.CTRL
flabel via3 18464 35376 24044 36196 0 FreeSans 1600 0 0 0 distortionUnit_2.VSS
flabel via3 18464 37316 24024 38056 0 FreeSans 1600 0 0 0 distortionUnit_2.VDD
flabel metal3 26744 37936 27064 39276 0 FreeSans 1600 0 0 0 distortionUnit_2.OUT
flabel metal3 17944 38416 18284 39136 0 FreeSans 1600 0 0 0 distortionUnit_2.IN
flabel metal2 25184 36756 25504 36976 0 FreeSans 1600 0 0 0 distortionUnit_2.tgate_1.IN
flabel metal2 25184 36276 25504 36496 0 FreeSans 1600 0 0 0 distortionUnit_2.tgate_1.OUT
flabel metal2 25184 37096 25724 37316 0 FreeSans 1600 0 0 0 distortionUnit_2.tgate_1.CTRLB
flabel metal2 25184 35936 25724 36156 0 FreeSans 1600 0 0 0 distortionUnit_2.tgate_1.CTRL
flabel metal1 26544 36756 26864 36976 0 FreeSans 1600 0 0 0 distortionUnit_2.tgate_1.VDD
flabel metal1 26544 36276 26864 36496 0 FreeSans 1600 0 0 0 distortionUnit_2.tgate_1.VSS
flabel metal2 25184 38216 25504 38436 0 FreeSans 1600 0 0 0 distortionUnit_2.tgate_0.IN
flabel metal2 25184 37736 25504 37956 0 FreeSans 1600 0 0 0 distortionUnit_2.tgate_0.OUT
flabel metal2 25184 38556 25724 38776 0 FreeSans 1600 0 0 0 distortionUnit_2.tgate_0.CTRLB
flabel metal2 25184 37396 25724 37616 0 FreeSans 1600 0 0 0 distortionUnit_2.tgate_0.CTRL
flabel metal1 26544 38216 26864 38436 0 FreeSans 1600 0 0 0 distortionUnit_2.tgate_0.VDD
flabel metal1 26544 37736 26864 37956 0 FreeSans 1600 0 0 0 distortionUnit_2.tgate_0.VSS
flabel metal1 26189 35010 26237 35036 0 FreeSans 200 0 0 0 distortionUnit_2.sky130_fd_sc_hd__tap_2_0.VGND
flabel metal1 26191 35557 26245 35579 0 FreeSans 200 0 0 0 distortionUnit_2.sky130_fd_sc_hd__tap_2_0.VPWR
flabel locali 26205 35455 26230 35480 0 FreeSans 250 0 0 0 distortionUnit_2.sky130_fd_sc_hd__tap_2_0.VPB
flabel locali 26290 35116 26325 35146 0 FreeSans 250 0 0 0 distortionUnit_2.sky130_fd_sc_hd__tap_2_0.VNB
flabel locali 26298 35449 26320 35478 0 FreeSans 250 0 0 0 distortionUnit_2.sky130_fd_sc_hd__tap_2_0.VPB
rlabel comment 26170 35024 26170 35024 4 distortionUnit_2.sky130_fd_sc_hd__tap_2_0.tap_2
rlabel metal1 26170 34976 26354 35072 1 distortionUnit_2.sky130_fd_sc_hd__tap_2_0.VGND
rlabel metal1 26170 35520 26354 35616 1 distortionUnit_2.sky130_fd_sc_hd__tap_2_0.VPWR
flabel locali 25555 35245 25589 35279 0 FreeSans 250 0 0 0 distortionUnit_2.sky130_fd_sc_hd__inv_8_0.A
flabel locali 25647 35245 25681 35279 0 FreeSans 250 0 0 0 distortionUnit_2.sky130_fd_sc_hd__inv_8_0.A
flabel locali 25739 35245 25773 35279 0 FreeSans 250 0 0 0 distortionUnit_2.sky130_fd_sc_hd__inv_8_0.A
flabel locali 25831 35245 25865 35279 0 FreeSans 250 0 0 0 distortionUnit_2.sky130_fd_sc_hd__inv_8_0.A
flabel locali 25923 35245 25957 35279 0 FreeSans 250 0 0 0 distortionUnit_2.sky130_fd_sc_hd__inv_8_0.A
flabel locali 26015 35245 26049 35279 0 FreeSans 250 0 0 0 distortionUnit_2.sky130_fd_sc_hd__inv_8_0.A
flabel locali 26107 35245 26141 35279 0 FreeSans 250 0 0 0 distortionUnit_2.sky130_fd_sc_hd__inv_8_0.Y
flabel locali 25371 35245 25405 35279 0 FreeSans 250 0 0 0 distortionUnit_2.sky130_fd_sc_hd__inv_8_0.Y
flabel pwell 25371 35007 25405 35041 0 FreeSans 200 0 0 0 distortionUnit_2.sky130_fd_sc_hd__inv_8_0.VNB
flabel nwell 25371 35551 25405 35585 0 FreeSans 200 0 0 0 distortionUnit_2.sky130_fd_sc_hd__inv_8_0.VPB
flabel metal1 25371 35007 25405 35041 0 FreeSans 200 0 0 0 distortionUnit_2.sky130_fd_sc_hd__inv_8_0.VGND
flabel metal1 25371 35551 25405 35585 0 FreeSans 200 0 0 0 distortionUnit_2.sky130_fd_sc_hd__inv_8_0.VPWR
rlabel comment 25342 35024 25342 35024 4 distortionUnit_2.sky130_fd_sc_hd__inv_8_0.inv_8
rlabel metal1 25342 34976 26170 35072 1 distortionUnit_2.sky130_fd_sc_hd__inv_8_0.VGND
rlabel metal1 25342 35520 26170 35616 1 distortionUnit_2.sky130_fd_sc_hd__inv_8_0.VPWR
flabel metal3 23024 36576 23414 36966 0 FreeSans 800 0 0 0 distortionUnit_2.myOpamp_0.INn
flabel metal3 20994 36866 22654 37116 0 FreeSans 800 0 0 0 distortionUnit_2.myOpamp_0.OUT
flabel metal3 20234 35966 23444 36216 0 FreeSans 800 0 0 0 distortionUnit_2.myOpamp_0.VSS
flabel metal3 20224 37266 23454 37536 0 FreeSans 800 0 0 0 distortionUnit_2.myOpamp_0.VDD
flabel metal3 20264 36866 20654 37176 0 FreeSans 800 0 0 0 distortionUnit_2.myOpamp_0.INp
flabel metal3 12532 18962 12892 19482 0 FreeSans 1600 0 0 0 distortionUnit_0.CTRL
flabel via3 5692 15582 11272 16402 0 FreeSans 1600 0 0 0 distortionUnit_0.VSS
flabel via3 5692 17522 11252 18262 0 FreeSans 1600 0 0 0 distortionUnit_0.VDD
flabel metal3 13972 18142 14292 19482 0 FreeSans 1600 0 0 0 distortionUnit_0.OUT
flabel metal3 5172 18622 5512 19342 0 FreeSans 1600 0 0 0 distortionUnit_0.IN
flabel metal2 12412 16962 12732 17182 0 FreeSans 1600 0 0 0 distortionUnit_0.tgate_1.IN
flabel metal2 12412 16482 12732 16702 0 FreeSans 1600 0 0 0 distortionUnit_0.tgate_1.OUT
flabel metal2 12412 17302 12952 17522 0 FreeSans 1600 0 0 0 distortionUnit_0.tgate_1.CTRLB
flabel metal2 12412 16142 12952 16362 0 FreeSans 1600 0 0 0 distortionUnit_0.tgate_1.CTRL
flabel metal1 13772 16962 14092 17182 0 FreeSans 1600 0 0 0 distortionUnit_0.tgate_1.VDD
flabel metal1 13772 16482 14092 16702 0 FreeSans 1600 0 0 0 distortionUnit_0.tgate_1.VSS
flabel metal2 12412 18422 12732 18642 0 FreeSans 1600 0 0 0 distortionUnit_0.tgate_0.IN
flabel metal2 12412 17942 12732 18162 0 FreeSans 1600 0 0 0 distortionUnit_0.tgate_0.OUT
flabel metal2 12412 18762 12952 18982 0 FreeSans 1600 0 0 0 distortionUnit_0.tgate_0.CTRLB
flabel metal2 12412 17602 12952 17822 0 FreeSans 1600 0 0 0 distortionUnit_0.tgate_0.CTRL
flabel metal1 13772 18422 14092 18642 0 FreeSans 1600 0 0 0 distortionUnit_0.tgate_0.VDD
flabel metal1 13772 17942 14092 18162 0 FreeSans 1600 0 0 0 distortionUnit_0.tgate_0.VSS
flabel metal1 13417 15216 13465 15242 0 FreeSans 200 0 0 0 distortionUnit_0.sky130_fd_sc_hd__tap_2_0.VGND
flabel metal1 13419 15763 13473 15785 0 FreeSans 200 0 0 0 distortionUnit_0.sky130_fd_sc_hd__tap_2_0.VPWR
flabel locali 13433 15661 13458 15686 0 FreeSans 250 0 0 0 distortionUnit_0.sky130_fd_sc_hd__tap_2_0.VPB
flabel locali 13518 15322 13553 15352 0 FreeSans 250 0 0 0 distortionUnit_0.sky130_fd_sc_hd__tap_2_0.VNB
flabel locali 13526 15655 13548 15684 0 FreeSans 250 0 0 0 distortionUnit_0.sky130_fd_sc_hd__tap_2_0.VPB
rlabel comment 13398 15230 13398 15230 4 distortionUnit_0.sky130_fd_sc_hd__tap_2_0.tap_2
rlabel metal1 13398 15182 13582 15278 1 distortionUnit_0.sky130_fd_sc_hd__tap_2_0.VGND
rlabel metal1 13398 15726 13582 15822 1 distortionUnit_0.sky130_fd_sc_hd__tap_2_0.VPWR
flabel locali 12783 15451 12817 15485 0 FreeSans 250 0 0 0 distortionUnit_0.sky130_fd_sc_hd__inv_8_0.A
flabel locali 12875 15451 12909 15485 0 FreeSans 250 0 0 0 distortionUnit_0.sky130_fd_sc_hd__inv_8_0.A
flabel locali 12967 15451 13001 15485 0 FreeSans 250 0 0 0 distortionUnit_0.sky130_fd_sc_hd__inv_8_0.A
flabel locali 13059 15451 13093 15485 0 FreeSans 250 0 0 0 distortionUnit_0.sky130_fd_sc_hd__inv_8_0.A
flabel locali 13151 15451 13185 15485 0 FreeSans 250 0 0 0 distortionUnit_0.sky130_fd_sc_hd__inv_8_0.A
flabel locali 13243 15451 13277 15485 0 FreeSans 250 0 0 0 distortionUnit_0.sky130_fd_sc_hd__inv_8_0.A
flabel locali 13335 15451 13369 15485 0 FreeSans 250 0 0 0 distortionUnit_0.sky130_fd_sc_hd__inv_8_0.Y
flabel locali 12599 15451 12633 15485 0 FreeSans 250 0 0 0 distortionUnit_0.sky130_fd_sc_hd__inv_8_0.Y
flabel pwell 12599 15213 12633 15247 0 FreeSans 200 0 0 0 distortionUnit_0.sky130_fd_sc_hd__inv_8_0.VNB
flabel nwell 12599 15757 12633 15791 0 FreeSans 200 0 0 0 distortionUnit_0.sky130_fd_sc_hd__inv_8_0.VPB
flabel metal1 12599 15213 12633 15247 0 FreeSans 200 0 0 0 distortionUnit_0.sky130_fd_sc_hd__inv_8_0.VGND
flabel metal1 12599 15757 12633 15791 0 FreeSans 200 0 0 0 distortionUnit_0.sky130_fd_sc_hd__inv_8_0.VPWR
rlabel comment 12570 15230 12570 15230 4 distortionUnit_0.sky130_fd_sc_hd__inv_8_0.inv_8
rlabel metal1 12570 15182 13398 15278 1 distortionUnit_0.sky130_fd_sc_hd__inv_8_0.VGND
rlabel metal1 12570 15726 13398 15822 1 distortionUnit_0.sky130_fd_sc_hd__inv_8_0.VPWR
flabel metal3 10252 16782 10642 17172 0 FreeSans 800 0 0 0 distortionUnit_0.myOpamp_0.INn
flabel metal3 8222 17072 9882 17322 0 FreeSans 800 0 0 0 distortionUnit_0.myOpamp_0.OUT
flabel metal3 7462 16172 10672 16422 0 FreeSans 800 0 0 0 distortionUnit_0.myOpamp_0.VSS
flabel metal3 7452 17472 10682 17742 0 FreeSans 800 0 0 0 distortionUnit_0.myOpamp_0.VDD
flabel metal3 7492 17072 7882 17382 0 FreeSans 800 0 0 0 distortionUnit_0.myOpamp_0.INp
flabel metal3 12516 38638 12876 39158 0 FreeSans 1600 0 0 0 bufferUnit_0.CTRL
flabel via3 5676 35258 11256 36078 0 FreeSans 1600 0 0 0 bufferUnit_0.VSS
flabel via3 5676 37198 11236 37938 0 FreeSans 1600 0 0 0 bufferUnit_0.VDD
flabel metal3 13956 37818 14276 39158 0 FreeSans 1600 0 0 0 bufferUnit_0.OUT
flabel metal3 5156 38298 5496 39018 0 FreeSans 1600 0 0 0 bufferUnit_0.IN
flabel metal2 12396 36638 12716 36858 0 FreeSans 1600 0 0 0 bufferUnit_0.tgate_1.IN
flabel metal2 12396 36158 12716 36378 0 FreeSans 1600 0 0 0 bufferUnit_0.tgate_1.OUT
flabel metal2 12396 36978 12936 37198 0 FreeSans 1600 0 0 0 bufferUnit_0.tgate_1.CTRLB
flabel metal2 12396 35818 12936 36038 0 FreeSans 1600 0 0 0 bufferUnit_0.tgate_1.CTRL
flabel metal1 13756 36638 14076 36858 0 FreeSans 1600 0 0 0 bufferUnit_0.tgate_1.VDD
flabel metal1 13756 36158 14076 36378 0 FreeSans 1600 0 0 0 bufferUnit_0.tgate_1.VSS
flabel metal2 12396 38098 12716 38318 0 FreeSans 1600 0 0 0 bufferUnit_0.tgate_0.IN
flabel metal2 12396 37618 12716 37838 0 FreeSans 1600 0 0 0 bufferUnit_0.tgate_0.OUT
flabel metal2 12396 38438 12936 38658 0 FreeSans 1600 0 0 0 bufferUnit_0.tgate_0.CTRLB
flabel metal2 12396 37278 12936 37498 0 FreeSans 1600 0 0 0 bufferUnit_0.tgate_0.CTRL
flabel metal1 13756 38098 14076 38318 0 FreeSans 1600 0 0 0 bufferUnit_0.tgate_0.VDD
flabel metal1 13756 37618 14076 37838 0 FreeSans 1600 0 0 0 bufferUnit_0.tgate_0.VSS
flabel metal1 13401 34892 13449 34918 0 FreeSans 200 0 0 0 bufferUnit_0.sky130_fd_sc_hd__tap_2_0.VGND
flabel metal1 13403 35439 13457 35461 0 FreeSans 200 0 0 0 bufferUnit_0.sky130_fd_sc_hd__tap_2_0.VPWR
flabel locali 13417 35337 13442 35362 0 FreeSans 250 0 0 0 bufferUnit_0.sky130_fd_sc_hd__tap_2_0.VPB
flabel locali 13502 34998 13537 35028 0 FreeSans 250 0 0 0 bufferUnit_0.sky130_fd_sc_hd__tap_2_0.VNB
flabel locali 13510 35331 13532 35360 0 FreeSans 250 0 0 0 bufferUnit_0.sky130_fd_sc_hd__tap_2_0.VPB
rlabel comment 13382 34906 13382 34906 4 bufferUnit_0.sky130_fd_sc_hd__tap_2_0.tap_2
rlabel metal1 13382 34858 13566 34954 1 bufferUnit_0.sky130_fd_sc_hd__tap_2_0.VGND
rlabel metal1 13382 35402 13566 35498 1 bufferUnit_0.sky130_fd_sc_hd__tap_2_0.VPWR
flabel locali 12767 35127 12801 35161 0 FreeSans 250 0 0 0 bufferUnit_0.sky130_fd_sc_hd__inv_8_0.A
flabel locali 12859 35127 12893 35161 0 FreeSans 250 0 0 0 bufferUnit_0.sky130_fd_sc_hd__inv_8_0.A
flabel locali 12951 35127 12985 35161 0 FreeSans 250 0 0 0 bufferUnit_0.sky130_fd_sc_hd__inv_8_0.A
flabel locali 13043 35127 13077 35161 0 FreeSans 250 0 0 0 bufferUnit_0.sky130_fd_sc_hd__inv_8_0.A
flabel locali 13135 35127 13169 35161 0 FreeSans 250 0 0 0 bufferUnit_0.sky130_fd_sc_hd__inv_8_0.A
flabel locali 13227 35127 13261 35161 0 FreeSans 250 0 0 0 bufferUnit_0.sky130_fd_sc_hd__inv_8_0.A
flabel locali 13319 35127 13353 35161 0 FreeSans 250 0 0 0 bufferUnit_0.sky130_fd_sc_hd__inv_8_0.Y
flabel locali 12583 35127 12617 35161 0 FreeSans 250 0 0 0 bufferUnit_0.sky130_fd_sc_hd__inv_8_0.Y
flabel pwell 12583 34889 12617 34923 0 FreeSans 200 0 0 0 bufferUnit_0.sky130_fd_sc_hd__inv_8_0.VNB
flabel nwell 12583 35433 12617 35467 0 FreeSans 200 0 0 0 bufferUnit_0.sky130_fd_sc_hd__inv_8_0.VPB
flabel metal1 12583 34889 12617 34923 0 FreeSans 200 0 0 0 bufferUnit_0.sky130_fd_sc_hd__inv_8_0.VGND
flabel metal1 12583 35433 12617 35467 0 FreeSans 200 0 0 0 bufferUnit_0.sky130_fd_sc_hd__inv_8_0.VPWR
rlabel comment 12554 34906 12554 34906 4 bufferUnit_0.sky130_fd_sc_hd__inv_8_0.inv_8
rlabel metal1 12554 34858 13382 34954 1 bufferUnit_0.sky130_fd_sc_hd__inv_8_0.VGND
rlabel metal1 12554 35402 13382 35498 1 bufferUnit_0.sky130_fd_sc_hd__inv_8_0.VPWR
flabel metal3 10236 36458 10626 36848 0 FreeSans 800 0 0 0 bufferUnit_0.myOpamp_0.INn
flabel metal3 8206 36748 9866 36998 0 FreeSans 800 0 0 0 bufferUnit_0.myOpamp_0.OUT
flabel metal3 7446 35848 10656 36098 0 FreeSans 800 0 0 0 bufferUnit_0.myOpamp_0.VSS
flabel metal3 7436 37148 10666 37418 0 FreeSans 800 0 0 0 bufferUnit_0.myOpamp_0.VDD
flabel metal3 7476 36748 7866 37058 0 FreeSans 800 0 0 0 bufferUnit_0.myOpamp_0.INp
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
