magic
tech sky130A
magscale 1 2
timestamp 1713223699
<< xpolycontact >>
rect -616 284 -546 716
rect -616 -716 -546 -284
rect -450 284 -380 716
rect -450 -716 -380 -284
rect -284 284 -214 716
rect -284 -716 -214 -284
rect -118 284 -48 716
rect -118 -716 -48 -284
rect 48 284 118 716
rect 48 -716 118 -284
rect 214 284 284 716
rect 214 -716 284 -284
rect 380 284 450 716
rect 380 -716 450 -284
rect 546 284 616 716
rect 546 -716 616 -284
<< xpolyres >>
rect -616 -284 -546 284
rect -450 -284 -380 284
rect -284 -284 -214 284
rect -118 -284 -48 284
rect 48 -284 118 284
rect 214 -284 284 284
rect 380 -284 450 284
rect 546 -284 616 284
<< viali >>
rect -600 301 -562 698
rect -434 301 -396 698
rect -268 301 -230 698
rect -102 301 -64 698
rect 64 301 102 698
rect 230 301 268 698
rect 396 301 434 698
rect 562 301 600 698
rect -600 -698 -562 -301
rect -434 -698 -396 -301
rect -268 -698 -230 -301
rect -102 -698 -64 -301
rect 64 -698 102 -301
rect 230 -698 268 -301
rect 396 -698 434 -301
rect 562 -698 600 -301
<< metal1 >>
rect -606 698 -556 710
rect -606 301 -600 698
rect -562 301 -556 698
rect -606 289 -556 301
rect -440 698 -390 710
rect -440 301 -434 698
rect -396 301 -390 698
rect -440 289 -390 301
rect -274 698 -224 710
rect -274 301 -268 698
rect -230 301 -224 698
rect -274 289 -224 301
rect -108 698 -58 710
rect -108 301 -102 698
rect -64 301 -58 698
rect -108 289 -58 301
rect 58 698 108 710
rect 58 301 64 698
rect 102 301 108 698
rect 58 289 108 301
rect 224 698 274 710
rect 224 301 230 698
rect 268 301 274 698
rect 224 289 274 301
rect 390 698 440 710
rect 390 301 396 698
rect 434 301 440 698
rect 390 289 440 301
rect 556 698 606 710
rect 556 301 562 698
rect 600 301 606 698
rect 556 289 606 301
rect -606 -301 -556 -289
rect -606 -698 -600 -301
rect -562 -698 -556 -301
rect -606 -710 -556 -698
rect -440 -301 -390 -289
rect -440 -698 -434 -301
rect -396 -698 -390 -301
rect -440 -710 -390 -698
rect -274 -301 -224 -289
rect -274 -698 -268 -301
rect -230 -698 -224 -301
rect -274 -710 -224 -698
rect -108 -301 -58 -289
rect -108 -698 -102 -301
rect -64 -698 -58 -301
rect -108 -710 -58 -698
rect 58 -301 108 -289
rect 58 -698 64 -301
rect 102 -698 108 -301
rect 58 -710 108 -698
rect 224 -301 274 -289
rect 224 -698 230 -301
rect 268 -698 274 -301
rect 224 -710 274 -698
rect 390 -301 440 -289
rect 390 -698 396 -301
rect 434 -698 440 -301
rect 390 -710 440 -698
rect 556 -301 606 -289
rect 556 -698 562 -301
rect 600 -698 606 -301
rect 556 -710 606 -698
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.35 l 3.0 m 1 nx 8 wmin 0.350 lmin 0.50 rho 2000 val 18.218k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 0 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
