magic
tech sky130A
magscale 1 2
timestamp 1713223699
<< nmos >>
rect -229 -19 -29 81
rect 29 -19 229 81
<< ndiff >>
rect -287 69 -229 81
rect -287 -7 -275 69
rect -241 -7 -229 69
rect -287 -19 -229 -7
rect -29 69 29 81
rect -29 -7 -17 69
rect 17 -7 29 69
rect -29 -19 29 -7
rect 229 69 287 81
rect 229 -7 241 69
rect 275 -7 287 69
rect 229 -19 287 -7
<< ndiffc >>
rect -275 -7 -241 69
rect -17 -7 17 69
rect 241 -7 275 69
<< poly >>
rect -229 81 -29 107
rect 29 81 229 107
rect -229 -57 -29 -19
rect -229 -91 -213 -57
rect -45 -91 -29 -57
rect -229 -107 -29 -91
rect 29 -57 229 -19
rect 29 -91 45 -57
rect 213 -91 229 -57
rect 29 -107 229 -91
<< polycont >>
rect -213 -91 -45 -57
rect 45 -91 213 -57
<< locali >>
rect -275 69 -241 85
rect -275 -23 -241 -7
rect -17 69 17 85
rect -17 -23 17 -7
rect 241 69 275 85
rect 241 -23 275 -7
rect -229 -91 -213 -57
rect -45 -91 -29 -57
rect 29 -91 45 -57
rect 213 -91 229 -57
<< viali >>
rect -275 -7 -241 69
rect -17 -7 17 69
rect 241 -7 275 69
rect -213 -91 -45 -57
rect 45 -91 213 -57
<< metal1 >>
rect -281 69 -235 81
rect -281 -7 -275 69
rect -241 -7 -235 69
rect -281 -19 -235 -7
rect -23 69 23 81
rect -23 -7 -17 69
rect 17 -7 23 69
rect -23 -19 23 -7
rect 235 69 281 81
rect 235 -7 241 69
rect 275 -7 281 69
rect 235 -19 281 -7
rect -225 -57 -33 -51
rect -225 -91 -213 -57
rect -45 -91 -33 -57
rect -225 -97 -33 -91
rect 33 -57 225 -51
rect 33 -91 45 -57
rect 213 -91 225 -57
rect 33 -97 225 -91
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.5 l 1 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
