magic
tech sky130A
magscale 1 2
timestamp 1713311859
<< nwell >>
rect 26 880 3252 1024
rect 26 849 3253 880
rect 25 835 3253 849
rect 25 512 312 835
rect 2985 511 3253 835
<< pwell >>
rect 20 -370 3250 -200
<< psubdiff >>
rect 70 -250 3200 -220
rect 70 -300 110 -250
rect 3160 -300 3200 -250
rect 70 -329 3200 -300
rect 70 -330 430 -329
rect 2840 -330 3200 -329
<< nsubdiff >>
rect 110 940 3200 980
rect 110 900 150 940
rect 3160 900 3200 940
rect 110 870 3200 900
<< psubdiffcont >>
rect 110 -300 3160 -250
<< nsubdiffcont >>
rect 150 900 3160 940
<< locali >>
rect -480 940 3210 980
rect -480 900 -420 940
rect 3160 900 3210 940
rect -480 860 3210 900
rect -480 -190 -40 -160
rect -480 -280 -460 -190
rect -60 -280 -40 -190
rect -480 -300 -40 -280
rect 70 -250 3210 -220
rect 70 -300 110 -250
rect 3160 -300 3210 -250
rect 70 -330 3210 -300
<< viali >>
rect -420 900 150 940
rect 150 900 3160 940
rect -460 -280 -60 -190
rect 110 -300 3160 -250
<< metal1 >>
rect -480 960 3210 980
rect -480 940 30 960
rect -480 900 -420 940
rect -480 880 30 900
rect 3190 880 3210 960
rect -480 860 3210 880
rect 70 570 130 860
rect 320 810 380 820
rect 280 690 430 810
rect 280 630 290 690
rect 400 630 430 690
rect 280 620 430 630
rect 540 620 670 860
rect 800 690 930 810
rect 800 630 810 690
rect 920 630 930 690
rect 800 620 930 630
rect 1060 620 1190 860
rect 1310 690 1440 820
rect 320 610 430 620
rect 70 530 320 570
rect 380 565 430 610
rect 1310 580 1320 690
rect 1430 580 1440 690
rect 1570 620 1700 860
rect 1830 700 1960 810
rect 1830 630 1840 700
rect 1950 630 1960 700
rect 1830 620 1960 630
rect 2090 620 2220 860
rect 2350 700 2480 820
rect 1310 565 1440 580
rect 2350 580 2360 700
rect 2470 580 2480 700
rect 2610 620 2740 860
rect 2860 700 2990 810
rect 2860 630 2870 700
rect 2980 630 2990 700
rect 2860 620 2990 630
rect 3170 580 3210 860
rect 2350 570 2480 580
rect 2360 565 2470 570
rect 378 531 2900 565
rect 380 530 430 531
rect 2960 530 3210 580
rect 660 480 770 490
rect 660 457 670 480
rect 378 423 670 457
rect 70 180 120 390
rect 280 370 410 380
rect 280 310 290 370
rect 400 310 410 370
rect 660 320 670 423
rect 760 457 770 480
rect 2730 480 2830 490
rect 760 423 2642 457
rect 760 320 770 423
rect 660 310 770 320
rect 800 370 930 380
rect 800 310 810 370
rect 920 310 930 370
rect 280 190 410 310
rect 540 260 670 280
rect 540 200 550 260
rect 660 200 670 260
rect 540 190 670 200
rect 800 190 930 310
rect 1060 260 1190 380
rect 1060 200 1070 260
rect 1180 200 1190 260
rect 1060 190 1190 200
rect 1310 370 1440 380
rect 1310 310 1320 370
rect 1430 310 1440 370
rect 1310 190 1440 310
rect 1580 260 1710 380
rect 1580 200 1590 260
rect 1700 200 1710 260
rect 1580 190 1710 200
rect 1830 370 1960 380
rect 1830 310 1840 370
rect 1950 310 1960 370
rect 1830 190 1960 310
rect 2090 260 2220 380
rect 2090 200 2100 260
rect 2210 200 2220 260
rect 2090 190 2220 200
rect 2350 370 2480 380
rect 2350 310 2360 370
rect 2470 310 2480 370
rect 2350 190 2480 310
rect 2730 330 2740 480
rect 2820 330 2830 480
rect 2730 300 2830 330
rect 2600 260 2730 270
rect 2600 200 2610 260
rect 2720 200 2730 260
rect 2600 190 2730 200
rect 70 150 140 180
rect 70 50 320 150
rect 2760 147 2830 300
rect 2860 370 2990 380
rect 2860 310 2870 370
rect 2980 310 2990 370
rect 2860 190 2990 310
rect 3160 180 3210 390
rect 3130 150 3210 180
rect 636 113 2900 147
rect 70 -47 840 50
rect 1520 40 1530 70
rect 890 10 1530 40
rect 1750 40 1760 70
rect 2950 50 3210 150
rect 1750 10 2390 40
rect 890 -19 2390 10
rect 1520 -30 1760 -19
rect -480 -170 -40 -160
rect -480 -290 -470 -170
rect -50 -290 -40 -170
rect -480 -300 -40 -290
rect 70 -220 884 -47
rect 1080 -125 1095 -47
rect 1150 -125 1170 -47
rect 1080 -135 1170 -125
rect 1310 -220 1450 -48
rect 1595 -140 1685 -30
rect 1830 -220 1970 -48
rect 2115 -125 2125 -48
rect 2180 -125 2190 -48
rect 2440 -50 3210 50
rect 2115 -135 2190 -125
rect 2390 -220 3210 -50
rect 70 -240 3210 -220
rect 70 -310 90 -240
rect 3190 -310 3210 -240
rect 70 -330 3210 -310
<< via1 >>
rect 30 940 3190 960
rect 30 900 3160 940
rect 3160 900 3190 940
rect 30 880 3190 900
rect 290 630 400 690
rect 810 630 920 690
rect 1320 580 1430 690
rect 1840 630 1950 700
rect 2360 580 2470 700
rect 2870 630 2980 700
rect 290 310 400 370
rect 670 320 760 480
rect 810 310 920 370
rect 550 200 660 260
rect 1070 200 1180 260
rect 1320 310 1430 370
rect 1590 200 1700 260
rect 1840 310 1950 370
rect 2100 200 2210 260
rect 2360 310 2470 370
rect 2740 330 2820 480
rect 2610 200 2720 260
rect 2870 310 2980 370
rect 1530 10 1750 70
rect -470 -190 -50 -170
rect -470 -280 -460 -190
rect -460 -280 -60 -190
rect -60 -280 -50 -190
rect -470 -290 -50 -280
rect 1095 -125 1150 -47
rect 2125 -125 2180 -48
rect 90 -250 3190 -240
rect 90 -300 110 -250
rect 110 -300 3160 -250
rect 3160 -300 3190 -250
rect 90 -310 3190 -300
<< metal2 >>
rect 10 1120 3260 1164
rect 10 850 20 1120
rect 3250 850 3260 1120
rect 10 840 3260 850
rect 280 690 410 700
rect 280 630 290 690
rect 400 630 410 690
rect 280 380 410 630
rect 280 310 290 380
rect 400 310 410 380
rect 280 300 410 310
rect 440 690 770 700
rect 440 470 450 690
rect 720 480 770 690
rect 440 320 670 470
rect 760 320 770 480
rect 440 300 770 320
rect 800 690 930 700
rect 800 620 810 690
rect 920 620 930 690
rect 800 370 930 620
rect 800 310 810 370
rect 920 310 930 370
rect 800 300 930 310
rect 1310 690 1440 710
rect 1310 580 1320 690
rect 1430 580 1440 690
rect 1310 380 1440 580
rect 1310 310 1320 380
rect 1430 310 1440 380
rect 1310 300 1440 310
rect 1830 700 1960 710
rect 1830 620 1840 700
rect 1950 620 1960 700
rect 1830 370 1960 620
rect 1830 310 1840 370
rect 1950 310 1960 370
rect 1830 300 1960 310
rect 2350 700 2480 710
rect 2350 580 2360 700
rect 2470 580 2480 700
rect 2350 380 2480 580
rect 2860 700 2990 710
rect 2860 620 2870 700
rect 2980 620 2990 700
rect 2350 310 2360 380
rect 2470 310 2480 380
rect 2530 490 2830 500
rect 2530 320 2550 490
rect 2820 320 2830 490
rect 2530 310 2830 320
rect 2860 370 2990 620
rect 2860 310 2870 370
rect 2980 310 2990 370
rect 2350 300 2480 310
rect 2860 300 2990 310
rect 530 260 2740 270
rect 530 200 550 260
rect 660 200 1070 260
rect 1180 200 1590 260
rect 1700 200 2100 260
rect 2210 200 2610 260
rect 2720 200 2740 260
rect 530 180 2740 200
rect -480 70 1780 110
rect -480 10 1530 70
rect 1750 10 1780 70
rect -480 0 1780 10
rect -480 -170 -40 0
rect 1850 -35 2210 180
rect 1060 -47 2210 -35
rect 1060 -125 1095 -47
rect 1150 -48 2210 -47
rect 1150 -125 2125 -48
rect 2180 -125 2210 -48
rect 1060 -140 2210 -125
rect -480 -290 -470 -170
rect -50 -290 -40 -170
rect -480 -300 -40 -290
rect 10 -450 30 -200
rect 3240 -450 3260 -200
rect 10 -568 3260 -450
<< via2 >>
rect 20 960 3250 1120
rect 20 880 30 960
rect 30 880 3190 960
rect 3190 880 3250 960
rect 20 850 3250 880
rect 290 370 400 380
rect 290 310 400 370
rect 450 480 720 690
rect 450 470 670 480
rect 670 470 720 480
rect 810 630 920 690
rect 810 620 920 630
rect 1320 370 1430 380
rect 1320 310 1430 370
rect 1840 630 1950 690
rect 1840 620 1950 630
rect 2870 630 2980 690
rect 2870 620 2980 630
rect 2360 370 2470 380
rect 2360 310 2470 370
rect 2550 480 2820 490
rect 2550 330 2740 480
rect 2740 330 2820 480
rect 2550 320 2820 330
rect 30 -240 3240 -200
rect 30 -310 90 -240
rect 90 -310 3190 -240
rect 3190 -310 3240 -240
rect 30 -450 3240 -310
<< metal3 >>
rect -1218 1120 3368 1164
rect -1218 850 20 1120
rect 3250 850 3368 1120
rect -1218 840 3368 850
rect 60 690 730 760
rect 60 470 450 690
rect 720 470 730 690
rect 60 450 730 470
rect 790 690 2990 700
rect 790 620 810 690
rect 920 620 1840 690
rect 1950 620 2870 690
rect 2980 620 2990 690
rect 790 610 2990 620
rect 790 450 2450 610
rect 2540 490 3210 550
rect 280 380 2480 390
rect 280 310 290 380
rect 400 310 1320 380
rect 1430 310 2360 380
rect 2470 310 2480 380
rect 280 300 2480 310
rect 820 140 2480 300
rect 2540 320 2550 490
rect 2820 320 3210 490
rect 2540 160 3210 320
rect -1218 -200 3368 -170
rect -1218 -450 30 -200
rect 3240 -450 3368 -200
rect -1218 -568 3368 -450
use sky130_fd_pr__nfet_01v8_7AMGGK  sky130_fd_pr__nfet_01v8_7AMGGK_0
timestamp 1713148837
transform 1 0 736 0 1 254
box -158 -157 158 157
use sky130_fd_pr__nfet_01v8_7AMGGK  sky130_fd_pr__nfet_01v8_7AMGGK_1
timestamp 1713148837
transform 1 0 2026 0 1 254
box -158 -157 158 157
use sky130_fd_pr__nfet_01v8_7AMGGK  sky130_fd_pr__nfet_01v8_7AMGGK_3
timestamp 1713148837
transform 1 0 2800 0 1 254
box -158 -157 158 157
use sky130_fd_pr__nfet_01v8_7AMGGK  sky130_fd_pr__nfet_01v8_7AMGGK_4
timestamp 1713148837
transform 1 0 1768 0 1 254
box -158 -157 158 157
use sky130_fd_pr__nfet_01v8_7AMGGK  sky130_fd_pr__nfet_01v8_7AMGGK_5
timestamp 1713148837
transform 1 0 994 0 1 254
box -158 -157 158 157
use sky130_fd_pr__nfet_01v8_7W2YM9  sky130_fd_pr__nfet_01v8_7W2YM9_0
timestamp 1713309734
transform 1 0 1639 0 1 -62
box -803 -99 803 99
use sky130_fd_pr__nfet_01v8_QFRGQ5  sky130_fd_pr__nfet_01v8_QFRGQ5_0
timestamp 1713148837
transform 1 0 478 0 1 316
box -158 -157 158 157
use sky130_fd_pr__nfet_01v8_QFRGQ5  sky130_fd_pr__nfet_01v8_QFRGQ5_1
timestamp 1713148837
transform 1 0 2284 0 1 316
box -158 -157 158 157
use sky130_fd_pr__nfet_01v8_QFRGQ5  sky130_fd_pr__nfet_01v8_QFRGQ5_2
timestamp 1713148837
transform 1 0 2542 0 1 316
box -158 -157 158 157
use sky130_fd_pr__nfet_01v8_QFRGQ5  sky130_fd_pr__nfet_01v8_QFRGQ5_3
timestamp 1713148837
transform 1 0 1252 0 1 316
box -158 -157 158 157
use sky130_fd_pr__nfet_01v8_QFRGQ5  sky130_fd_pr__nfet_01v8_QFRGQ5_5
timestamp 1713148837
transform 1 0 1510 0 1 316
box -158 -157 158 157
use sky130_fd_pr__pfet_01v8_PE7Z8M  sky130_fd_pr__pfet_01v8_PE7Z8M_0
timestamp 1713148837
transform 1 0 1639 0 1 676
box -1355 -164 1355 198
<< labels >>
flabel metal3 2820 160 3210 550 0 FreeSans 800 0 0 0 INn
port 5 nsew
flabel metal3 790 450 2450 700 0 FreeSans 800 0 0 0 OUT
port 1 nsew
flabel metal3 30 -450 3240 -200 0 FreeSans 800 0 0 0 VSS
port 2 nsew
flabel metal3 20 850 3250 1120 0 FreeSans 800 0 0 0 VDD
port 3 nsew
flabel metal3 60 450 450 760 0 FreeSans 800 0 0 0 INp
port 4 nsew
flabel metal2 -480 -170 -40 110 0 FreeSans 1600 0 0 0 R
port 6 nsew
<< end >>
