magic
tech sky130A
magscale 1 2
timestamp 1713148837
<< nwell >>
rect -1355 -164 1355 198
<< pmos >>
rect -1261 -64 -1061 136
rect -1003 -64 -803 136
rect -745 -64 -545 136
rect -487 -64 -287 136
rect -229 -64 -29 136
rect 29 -64 229 136
rect 287 -64 487 136
rect 545 -64 745 136
rect 803 -64 1003 136
rect 1061 -64 1261 136
<< pdiff >>
rect -1319 124 -1261 136
rect -1319 -52 -1307 124
rect -1273 -52 -1261 124
rect -1319 -64 -1261 -52
rect -1061 124 -1003 136
rect -1061 -52 -1049 124
rect -1015 -52 -1003 124
rect -1061 -64 -1003 -52
rect -803 124 -745 136
rect -803 -52 -791 124
rect -757 -52 -745 124
rect -803 -64 -745 -52
rect -545 124 -487 136
rect -545 -52 -533 124
rect -499 -52 -487 124
rect -545 -64 -487 -52
rect -287 124 -229 136
rect -287 -52 -275 124
rect -241 -52 -229 124
rect -287 -64 -229 -52
rect -29 124 29 136
rect -29 -52 -17 124
rect 17 -52 29 124
rect -29 -64 29 -52
rect 229 124 287 136
rect 229 -52 241 124
rect 275 -52 287 124
rect 229 -64 287 -52
rect 487 124 545 136
rect 487 -52 499 124
rect 533 -52 545 124
rect 487 -64 545 -52
rect 745 124 803 136
rect 745 -52 757 124
rect 791 -52 803 124
rect 745 -64 803 -52
rect 1003 124 1061 136
rect 1003 -52 1015 124
rect 1049 -52 1061 124
rect 1003 -64 1061 -52
rect 1261 124 1319 136
rect 1261 -52 1273 124
rect 1307 -52 1319 124
rect 1261 -64 1319 -52
<< pdiffc >>
rect -1307 -52 -1273 124
rect -1049 -52 -1015 124
rect -791 -52 -757 124
rect -533 -52 -499 124
rect -275 -52 -241 124
rect -17 -52 17 124
rect 241 -52 275 124
rect 499 -52 533 124
rect 757 -52 791 124
rect 1015 -52 1049 124
rect 1273 -52 1307 124
<< poly >>
rect -1261 136 -1061 162
rect -1003 136 -803 162
rect -745 136 -545 162
rect -487 136 -287 162
rect -229 136 -29 162
rect 29 136 229 162
rect 287 136 487 162
rect 545 136 745 162
rect 803 136 1003 162
rect 1061 136 1261 162
rect -1261 -111 -1061 -64
rect -1261 -145 -1245 -111
rect -1077 -145 -1061 -111
rect -1261 -161 -1061 -145
rect -1003 -111 -803 -64
rect -1003 -145 -987 -111
rect -819 -145 -803 -111
rect -1003 -161 -803 -145
rect -745 -111 -545 -64
rect -745 -145 -729 -111
rect -561 -145 -545 -111
rect -745 -161 -545 -145
rect -487 -111 -287 -64
rect -487 -145 -471 -111
rect -303 -145 -287 -111
rect -487 -161 -287 -145
rect -229 -111 -29 -64
rect -229 -145 -213 -111
rect -45 -145 -29 -111
rect -229 -161 -29 -145
rect 29 -111 229 -64
rect 29 -145 45 -111
rect 213 -145 229 -111
rect 29 -161 229 -145
rect 287 -111 487 -64
rect 287 -145 303 -111
rect 471 -145 487 -111
rect 287 -161 487 -145
rect 545 -111 745 -64
rect 545 -145 561 -111
rect 729 -145 745 -111
rect 545 -161 745 -145
rect 803 -111 1003 -64
rect 803 -145 819 -111
rect 987 -145 1003 -111
rect 803 -161 1003 -145
rect 1061 -111 1261 -64
rect 1061 -145 1077 -111
rect 1245 -145 1261 -111
rect 1061 -161 1261 -145
<< polycont >>
rect -1245 -145 -1077 -111
rect -987 -145 -819 -111
rect -729 -145 -561 -111
rect -471 -145 -303 -111
rect -213 -145 -45 -111
rect 45 -145 213 -111
rect 303 -145 471 -111
rect 561 -145 729 -111
rect 819 -145 987 -111
rect 1077 -145 1245 -111
<< locali >>
rect -1307 124 -1273 140
rect -1307 -68 -1273 -52
rect -1049 124 -1015 140
rect -1049 -68 -1015 -52
rect -791 124 -757 140
rect -791 -68 -757 -52
rect -533 124 -499 140
rect -533 -68 -499 -52
rect -275 124 -241 140
rect -275 -68 -241 -52
rect -17 124 17 140
rect -17 -68 17 -52
rect 241 124 275 140
rect 241 -68 275 -52
rect 499 124 533 140
rect 499 -68 533 -52
rect 757 124 791 140
rect 757 -68 791 -52
rect 1015 124 1049 140
rect 1015 -68 1049 -52
rect 1273 124 1307 140
rect 1273 -68 1307 -52
rect -1261 -145 -1245 -111
rect -1077 -145 -1061 -111
rect -1003 -145 -987 -111
rect -819 -145 -803 -111
rect -745 -145 -729 -111
rect -561 -145 -545 -111
rect -487 -145 -471 -111
rect -303 -145 -287 -111
rect -229 -145 -213 -111
rect -45 -145 -29 -111
rect 29 -145 45 -111
rect 213 -145 229 -111
rect 287 -145 303 -111
rect 471 -145 487 -111
rect 545 -145 561 -111
rect 729 -145 745 -111
rect 803 -145 819 -111
rect 987 -145 1003 -111
rect 1061 -145 1077 -111
rect 1245 -145 1261 -111
<< viali >>
rect -1307 -52 -1273 124
rect -1049 -52 -1015 124
rect -791 -52 -757 124
rect -533 -52 -499 124
rect -275 -52 -241 124
rect -17 -52 17 124
rect 241 -52 275 124
rect 499 -52 533 124
rect 757 -52 791 124
rect 1015 -52 1049 124
rect 1273 -52 1307 124
rect -1245 -145 -1077 -111
rect -987 -145 -819 -111
rect -729 -145 -561 -111
rect -471 -145 -303 -111
rect -213 -145 -45 -111
rect 45 -145 213 -111
rect 303 -145 471 -111
rect 561 -145 729 -111
rect 819 -145 987 -111
rect 1077 -145 1245 -111
<< metal1 >>
rect -1313 124 -1267 136
rect -1313 -52 -1307 124
rect -1273 -52 -1267 124
rect -1313 -64 -1267 -52
rect -1055 124 -1009 136
rect -1055 -52 -1049 124
rect -1015 -52 -1009 124
rect -1055 -64 -1009 -52
rect -797 124 -751 136
rect -797 -52 -791 124
rect -757 -52 -751 124
rect -797 -64 -751 -52
rect -539 124 -493 136
rect -539 -52 -533 124
rect -499 -52 -493 124
rect -539 -64 -493 -52
rect -281 124 -235 136
rect -281 -52 -275 124
rect -241 -52 -235 124
rect -281 -64 -235 -52
rect -23 124 23 136
rect -23 -52 -17 124
rect 17 -52 23 124
rect -23 -64 23 -52
rect 235 124 281 136
rect 235 -52 241 124
rect 275 -52 281 124
rect 235 -64 281 -52
rect 493 124 539 136
rect 493 -52 499 124
rect 533 -52 539 124
rect 493 -64 539 -52
rect 751 124 797 136
rect 751 -52 757 124
rect 791 -52 797 124
rect 751 -64 797 -52
rect 1009 124 1055 136
rect 1009 -52 1015 124
rect 1049 -52 1055 124
rect 1009 -64 1055 -52
rect 1267 124 1313 136
rect 1267 -52 1273 124
rect 1307 -52 1313 124
rect 1267 -64 1313 -52
rect -1257 -111 -1065 -105
rect -1257 -145 -1245 -111
rect -1077 -145 -1065 -111
rect -1257 -151 -1065 -145
rect -999 -111 -807 -105
rect -999 -145 -987 -111
rect -819 -145 -807 -111
rect -999 -151 -807 -145
rect -741 -111 -549 -105
rect -741 -145 -729 -111
rect -561 -145 -549 -111
rect -741 -151 -549 -145
rect -483 -111 -291 -105
rect -483 -145 -471 -111
rect -303 -145 -291 -111
rect -483 -151 -291 -145
rect -225 -111 -33 -105
rect -225 -145 -213 -111
rect -45 -145 -33 -111
rect -225 -151 -33 -145
rect 33 -111 225 -105
rect 33 -145 45 -111
rect 213 -145 225 -111
rect 33 -151 225 -145
rect 291 -111 483 -105
rect 291 -145 303 -111
rect 471 -145 483 -111
rect 291 -151 483 -145
rect 549 -111 741 -105
rect 549 -145 561 -111
rect 729 -145 741 -111
rect 549 -151 741 -145
rect 807 -111 999 -105
rect 807 -145 819 -111
rect 987 -145 999 -111
rect 807 -151 999 -145
rect 1065 -111 1257 -105
rect 1065 -145 1077 -111
rect 1245 -145 1257 -111
rect 1065 -151 1257 -145
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 1 m 1 nf 10 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
