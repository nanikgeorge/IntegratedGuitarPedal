magic
tech sky130A
magscale 1 2
timestamp 1713492510
<< locali >>
rect 5620 2720 5780 2740
rect 5620 2320 5640 2720
rect 5760 2320 5780 2720
rect 5620 2300 5780 2320
rect 5420 1180 5560 1200
rect 5420 740 5440 1180
rect 5540 740 5560 1180
rect 5420 720 5560 740
rect 3520 180 4680 200
rect 3520 100 3540 180
rect 4660 100 4680 180
rect 3520 80 4680 100
rect 5360 -220 5560 100
<< viali >>
rect 5640 2320 5760 2720
rect 5440 740 5540 1180
rect 6702 250 7190 284
rect 7314 184 7362 348
rect 3540 100 4660 180
<< metal1 >>
rect 7840 3420 8680 3480
rect 7840 3200 8560 3420
rect 8640 3200 8680 3420
rect 7840 3180 8680 3200
rect 7840 2960 8680 3000
rect 5580 2780 5840 2800
rect 5580 2300 5600 2780
rect 5820 2300 5840 2780
rect 7840 2740 8380 2960
rect 8460 2740 8680 2960
rect 7840 2700 8680 2740
rect 5580 2280 5840 2300
rect 7840 1960 8680 2020
rect 7840 1740 8560 1960
rect 8640 1740 8680 1960
rect 7840 1720 8680 1740
rect 7840 1500 8680 1540
rect 7840 1280 8380 1500
rect 8460 1280 8680 1500
rect 7840 1240 8680 1280
rect 5420 1180 5560 1200
rect 5420 740 5440 1180
rect 5540 740 5560 1180
rect 5420 720 5560 740
rect 6200 360 7200 380
rect 5600 320 5800 340
rect 3520 198 4680 200
rect 3516 180 4680 198
rect 3516 100 3540 180
rect 4660 100 4680 180
rect 3516 80 4680 100
rect 3516 -114 4104 80
rect 5600 60 5620 320
rect 4820 40 5620 60
rect 4820 -140 4840 40
rect 5780 -140 5800 320
rect 6200 180 6220 360
rect 6400 284 7200 360
rect 6400 250 6702 284
rect 7190 250 7200 284
rect 6400 180 7200 250
rect 6200 160 7200 180
rect 7300 360 7700 380
rect 7300 348 7500 360
rect 7300 184 7314 348
rect 7362 184 7500 348
rect 7300 180 7500 184
rect 7680 180 7700 360
rect 7300 160 7700 180
rect 4820 -160 5800 -140
<< via1 >>
rect 8560 3200 8640 3420
rect 5600 2720 5820 2780
rect 5600 2320 5640 2720
rect 5640 2320 5760 2720
rect 5760 2320 5820 2720
rect 5600 2300 5820 2320
rect 8380 2740 8460 2960
rect 8560 1740 8640 1960
rect 8380 1280 8460 1500
rect 5440 740 5540 1180
rect 6580 540 7540 600
rect 3540 100 4660 180
rect 5620 40 5780 320
rect 4840 -140 5780 40
rect 6220 180 6400 360
rect 7500 180 7680 360
rect 6580 0 7560 60
<< metal2 >>
rect -840 3420 6420 3440
rect -840 3240 -820 3420
rect -520 3240 6420 3420
rect -840 3220 6420 3240
rect 8540 3420 8660 3440
rect 8540 3200 8560 3420
rect 8640 3200 8660 3420
rect 8540 3180 8660 3200
rect 8360 2960 8480 2980
rect 7620 2940 8280 2960
rect 5580 2780 5840 2800
rect 5580 2300 5600 2780
rect 5820 2300 5840 2780
rect 7620 2760 7980 2940
rect 8260 2760 8280 2940
rect 7620 2740 8280 2760
rect 8360 2740 8380 2960
rect 8460 2740 8480 2960
rect 8360 2720 8480 2740
rect 5580 2280 5840 2300
rect 6400 2600 7780 2620
rect 6400 2120 7500 2600
rect 7680 2120 7780 2600
rect 6400 2100 7780 2120
rect 5940 1960 6540 1980
rect 5940 1780 5960 1960
rect 6160 1780 6540 1960
rect 5940 1760 6540 1780
rect 8540 1960 8660 1980
rect 8540 1740 8560 1960
rect 8640 1740 8660 1960
rect 8540 1720 8660 1740
rect 8360 1500 8480 1520
rect 7600 1480 8280 1500
rect 7600 1300 7980 1480
rect 8260 1300 8280 1480
rect 7600 1280 8280 1300
rect 8360 1280 8380 1500
rect 8460 1280 8480 1500
rect 8360 1260 8480 1280
rect 4660 1180 5580 1220
rect 4660 880 5440 1180
rect 3520 740 5440 880
rect 5540 740 5580 1180
rect 3520 700 5580 740
rect 6460 700 7580 720
rect 3520 180 4680 700
rect 6460 600 6980 700
rect 7360 600 7580 700
rect 6460 540 6580 600
rect 7540 540 7580 600
rect 6460 520 7580 540
rect 6200 360 6420 380
rect 3520 100 3540 180
rect 4660 100 4680 180
rect 3520 60 4680 100
rect 5600 320 5800 340
rect 5600 60 5620 320
rect 4820 40 5620 60
rect 4820 -140 4840 40
rect 5780 -140 5800 320
rect 6200 180 6220 360
rect 6400 180 6420 360
rect 6200 160 6420 180
rect 7480 360 7700 380
rect 7480 180 7500 360
rect 7680 180 7700 360
rect 7480 160 7700 180
rect 6460 60 7580 80
rect 6460 -100 6540 60
rect 7560 0 7580 60
rect 6860 -100 7580 0
rect 6460 -120 7580 -100
rect 4820 -160 5800 -140
<< via2 >>
rect 6540 3580 6860 3760
rect -820 3240 -520 3420
rect 8560 3200 8640 3420
rect 5600 2300 5820 2780
rect 7980 2760 8260 2940
rect 8380 2740 8460 2960
rect 7500 2120 7680 2600
rect 5960 1780 6160 1960
rect 8560 1740 8640 1960
rect 7980 1300 8260 1480
rect 8380 1280 8460 1500
rect 6460 960 6860 1140
rect 6980 600 7360 700
rect 6980 540 7360 600
rect 5620 40 5780 320
rect 4840 -140 5780 40
rect 6220 180 6400 360
rect 7500 180 7680 360
rect 6540 0 6580 60
rect 6580 0 6860 60
rect 6540 -100 6860 0
<< metal3 >>
rect -840 3420 -500 4140
rect -840 3240 -820 3420
rect -520 3240 -500 3420
rect -840 2180 -500 3240
rect 6520 3760 6880 4280
rect 6520 3580 6540 3760
rect 6860 3580 6880 3760
rect 5580 2780 5840 2800
rect 5580 2300 5600 2780
rect 5820 2300 5840 2780
rect 5580 2240 5840 2300
rect -840 1880 1860 2180
rect 5580 2140 6180 2240
rect 4040 2040 6180 2140
rect 5940 1960 6180 2040
rect 4240 1580 5800 1960
rect 5940 1780 5960 1960
rect 6160 1780 6180 1960
rect 5940 1760 6180 1780
rect 5600 320 5800 1580
rect 6520 1200 6880 3580
rect 5600 60 5620 320
rect 4820 40 5620 60
rect 4820 -140 4840 40
rect 5780 -140 5800 320
rect 6200 1140 6880 1200
rect 6200 960 6460 1140
rect 6860 960 6880 1140
rect 6200 880 6880 960
rect 6960 3100 7380 3120
rect 6960 2280 6980 3100
rect 7360 2280 7380 3100
rect 7960 2940 8280 4280
rect 8540 3420 8660 3440
rect 8540 3200 8560 3420
rect 8640 3200 8660 3420
rect 8540 3100 8660 3200
rect 7960 2760 7980 2940
rect 8260 2760 8280 2940
rect 6200 360 6420 880
rect 6200 180 6220 360
rect 6400 180 6420 360
rect 6200 160 6420 180
rect 6520 700 6880 720
rect 6520 340 6540 700
rect 6860 340 6880 700
rect 6960 700 7380 2280
rect 6960 540 6980 700
rect 7360 540 7380 700
rect 6960 520 7380 540
rect 7480 2600 7700 2620
rect 7480 2120 7500 2600
rect 7680 2120 7700 2600
rect 6520 60 6880 340
rect 7480 360 7700 2120
rect 7960 1480 8280 2760
rect 7960 1300 7980 1480
rect 8260 1300 8280 1480
rect 7960 1280 8280 1300
rect 8360 2960 8480 2980
rect 8360 2740 8380 2960
rect 8460 2740 8480 2960
rect 8360 1500 8480 2740
rect 8540 2280 8560 3100
rect 8640 2280 8660 3100
rect 8540 1960 8660 2280
rect 8540 1740 8560 1960
rect 8640 1740 8660 1960
rect 8540 1720 8660 1740
rect 8360 1280 8380 1500
rect 8460 1280 8480 1500
rect 7480 180 7500 360
rect 7680 180 7700 360
rect 8360 1240 8480 1280
rect 8360 340 8380 1240
rect 8460 340 8480 1240
rect 8360 320 8480 340
rect 7480 160 7700 180
rect 6520 -100 6540 60
rect 6860 -100 6880 60
rect 6520 -120 6880 -100
rect 4820 -160 5800 -140
<< via3 >>
rect -320 2320 5240 3060
rect -320 380 5260 1200
rect 6980 2280 7360 3100
rect 6540 340 6860 700
rect 8560 2280 8640 3100
rect 8380 340 8460 1240
<< metal4 >>
rect -380 3100 9200 3120
rect -380 3060 6980 3100
rect -380 2320 -320 3060
rect 5240 2320 6980 3060
rect -380 2280 6980 2320
rect 7360 2280 8560 3100
rect 8640 2280 9200 3100
rect -380 2260 9200 2280
rect -380 1240 9200 1260
rect -380 1200 8380 1240
rect -380 380 -320 1200
rect 5260 700 8380 1200
rect 5260 380 6540 700
rect -380 340 6540 380
rect 6860 340 8380 700
rect 8460 340 9200 1240
rect -380 320 9200 340
use inverter  inverter_0
timestamp 1713492510
transform 1 0 6613 0 1 -514
box 178 804 568 867
use myOpamp  myOpamp_0
timestamp 1713445313
transform 1 0 1420 0 1 1420
box -1800 -1100 3900 1700
use sky130_fd_pr__res_xhigh_po_0p69_FXQCTT  sky130_fd_pr__res_xhigh_po_0p69_FXQCTT_0
timestamp 1713488381
transform 0 -1 4442 1 0 -25
box -235 -982 235 982
use sky130_fd_pr__res_xhigh_po_0p69_WUKAVR  sky130_fd_pr__res_xhigh_po_0p69_WUKAVR_0
timestamp 1713488381
transform 1 0 5695 0 1 1322
box -235 -1582 235 1582
use sky130_fd_sc_hd__inv_8  sky130_fd_sc_hd__inv_8_0 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6558 0 1 28
box -38 -48 866 592
use sky130_fd_sc_hd__tap_2  sky130_fd_sc_hd__tap_2_0 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7386 0 1 28
box -38 -48 222 592
use tgate  tgate_0
timestamp 1713408040
transform 1 0 6780 0 1 2580
box -380 -180 1300 1200
use tgate  tgate_1
timestamp 1713408040
transform 1 0 6780 0 1 1120
box -380 -180 1300 1200
<< labels >>
flabel metal3 6520 3760 6880 4280 0 FreeSans 1600 0 0 0 CTRL
port 2 nsew
flabel via3 -320 380 5260 1200 0 FreeSans 1600 0 0 0 VSS
port 5 nsew
flabel via3 -320 2320 5240 3060 0 FreeSans 1600 0 0 0 VDD
port 4 nsew
flabel metal3 7960 2940 8280 4280 0 FreeSans 1600 0 0 0 OUT
port 3 nsew
flabel metal3 -840 3420 -500 4140 0 FreeSans 1600 0 0 0 IN
port 1 nsew
<< end >>
