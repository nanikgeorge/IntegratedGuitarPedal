* NGSPICE file created from guitflat7.ext - technology: sky130A

.subckt tt_um_guitar_pedal ua[0] ua[1] ui_in[0] VPWR ui_in[1] VGND ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7]
X0 VGND.t17 ui_in[4].t0 distortionUnit_5.tgate_1.CTRLB VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_20524_36601# a_20524_36601# VPWR.t76 VPWR.t75 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2 VGND.t378 VGND.t376 VGND.t378 VGND.t377 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X3 distortionUnit_0.tgate_1.CTRLB ui_in[6].t0 VPWR.t281 distortionUnit_0.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR.t276 VPWR.t274 distortionUnit_0.tgate_1.IN VPWR.t275 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X5 a_7876_23853# VGND.t374 VGND.t375 VGND.t301 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X6 VGND.t373 VGND.t372 VGND.t373 VGND.t42 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X7 VPWR.t132 a_7752_16807# a_7752_16807# VPWR.t131 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X8 distortionUnit_4.IN ui_in[3].t0 distortionUnit_5.IN.t5 VPWR.t278 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X9 ua[1].t3 ui_in[7].t0 distortionUnit_7.IN VPWR.t90 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X10 distortionUnit_6.IN ui_in[4].t1 distortionUnit_5.tgate_1.IN VGND.t15 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X11 a_7752_16807# distortionUnit_6.OUT a_8010_16807# VGND.t101 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X12 distortionUnit_4.tgate_1.IN distortionUnit_4.myOpamp_0.INn a_20746_30481# VGND.t157 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X13 VPWR.t184 a_20934_16677# distortionUnit_7.tgate_1.IN VPWR.t183 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X14 ua[1].t7 distortionUnit_7.tgate_1.CTRLB distortionUnit_7.IN VGND.t458 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X15 VPWR.t228 ui_in[0].t0 bufferUnit_0.tgate_1.CTRLB bufferUnit_0.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 VGND.t371 VGND.t369 VGND.t371 VGND.t370 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X17 distortionUnit_7.tgate_1.IN distortionUnit_7.myOpamp_0.INn a_21192_16677# VGND.t200 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X18 a_7752_16807# distortionUnit_6.OUT a_8010_16807# VGND.t99 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X19 VPWR.t99 ui_in[2].t0 distortionUnit_3.tgate_1.CTRLB distortionUnit_3.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 bufferUnit_0.tgate_1.IN bufferUnit_0.tgate_1.CTRLB bufferUnit_0.OUT VPWR.t79 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X21 VPWR.t282 ui_in[6].t1 distortionUnit_0.tgate_1.CTRLB distortionUnit_0.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X22 distortionUnit_6.tgate_1.CTRLB ui_in[5].t0 VPWR.t112 distortionUnit_6.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 VGND.t447 a_19680_36146# a_20782_36601# VGND.t446 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X24 distortionUnit_0.tgate_1.IN a_7752_16807# VPWR.t130 VPWR.t129 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X25 VGND.t450 ui_in[3].t1 distortionUnit_4.tgate_1.CTRLB VGND.t449 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 a_7994_36483# ua[0].t4 a_7736_36483# VGND.t293 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X27 distortionUnit_4.tgate_1.CTRLB ui_in[3].t2 VGND.t452 VGND.t451 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X28 a_20782_36601# distortionUnit_2.myOpamp_0.INn distortionUnit_2.tgate_1.IN VGND.t408 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X29 VPWR.t283 ui_in[6].t2 distortionUnit_0.tgate_1.CTRLB distortionUnit_0.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 VGND.t162 a_19644_30026# a_20746_30481# VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X31 distortionUnit_7.IN ui_in[6].t3 distortionUnit_6.OUT VPWR.t284 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X32 distortionUnit_7.IN distortionUnit_7.tgate_1.CTRLB ua[1].t6 VGND.t457 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X33 a_7752_16807# VPWR.t271 VPWR.t273 VPWR.t272 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X34 distortionUnit_6.tgate_1.IN ui_in[5].t1 distortionUnit_6.OUT VGND.t140 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X35 distortionUnit_3.tgate_1.CTRLB ui_in[2].t1 VPWR.t100 distortionUnit_3.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X36 a_7876_23853# a_7876_23853# VPWR.t32 VPWR.t31 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X37 VPWR.t270 VPWR.t268 distortionUnit_7.tgate_1.IN VPWR.t269 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X38 a_8010_16807# distortionUnit_0.myOpamp_0.INn distortionUnit_0.tgate_1.IN VGND.t97 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X39 a_20746_30481# distortionUnit_4.IN a_20488_30481# VGND.t44 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X40 VGND.t468 a_6912_30102# a_8014_30557# VGND.t75 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X41 VPWR.t311 a_7756_30557# a_7756_30557# VPWR.t310 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X42 a_7994_36483# a_6892_36028# VGND.t419 VGND.t418 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X43 VGND.t399 a_20090_16222# a_21192_16677# VGND.t203 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X44 distortionUnit_3.tgate_1.CTRLB ui_in[2].t2 VPWR.t101 distortionUnit_3.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X45 VGND.t368 VGND.t367 distortionUnit_3.tgate_1.IN VGND.t288 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X46 distortionUnit_5.tgate_1.CTRLB ui_in[4].t2 VGND.t14 VGND.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X47 distortionUnit_6.tgate_1.IN distortionUnit_6.myOpamp_0.INn a_20842_23723# VGND.t285 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X48 VPWR.t267 VPWR.t265 distortionUnit_2.tgate_1.IN VPWR.t266 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X49 distortionUnit_0.tgate_1.CTRLB ui_in[6].t4 VPWR.t42 distortionUnit_0.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X50 VGND distortionUnit_5.myOpamp_0.INn VGND.t88 sky130_fd_pr__res_xhigh_po_0p69 l=4
X51 a_8134_23853# distortionUnit_5.myOpamp_0.INn distortionUnit_5.tgate_1.IN VGND.t95 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X52 a_20782_36601# a_19680_36146# VGND.t445 VGND.t407 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X53 a_8014_30557# distortionUnit_3.IN a_7756_30557# VGND.t77 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X54 VPWR a_19680_36146# VGND sky130_fd_pr__res_xhigh_po_0p35 l=26.11
X55 distortionUnit_4.tgate_1.CTRLB ui_in[3].t3 VGND.t454 VGND.t453 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X56 VGND.t366 VGND.t365 VGND.t366 VGND.t332 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X57 VPWR.t277 a_19740_23268# VGND.t448 sky130_fd_pr__res_xhigh_po_0p35 l=0.16
X58 a_7736_36483# ua[0].t5 a_7994_36483# VGND.t413 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X59 distortionUnit_5.tgate_1.CTRLB ui_in[4].t3 VGND.t12 VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X60 distortionUnit_6.OUT distortionUnit_0.tgate_1.CTRLB distortionUnit_7.IN VGND.t393 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X61 bufferUnit_0.OUT ui_in[1].t0 distortionUnit_3.IN VPWR.t287 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X62 a_6908_16352# a_6908_16352# VGND.t108 VGND.t107 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X63 VGND.t173 ui_in[0].t1 bufferUnit_0.tgate_1.CTRLB VGND.t172 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X64 distortionUnit_7.tgate_1.IN a_20934_16677# VPWR.t182 VPWR.t181 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X65 VGND.t460 ui_in[1].t1 distortionUnit_2.tgate_1.CTRLB VGND.t459 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X66 distortionUnit_4.tgate_1.IN a_20488_30481# VPWR.t156 VPWR.t155 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X67 distortionUnit_6.tgate_1.IN a_20584_23723# VPWR.t205 VPWR.t204 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X68 distortionUnit_2.tgate_1.CTRLB ui_in[1].t2 VGND.t462 VGND.t461 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X69 a_21192_16677# a_20090_16222# VGND.t398 VGND.t199 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X70 distortionUnit_7.tgate_1.IN a_20934_16677# VPWR.t180 VPWR.t179 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X71 VPWR.t30 a_7876_23853# distortionUnit_5.tgate_1.IN VPWR.t29 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X72 distortionUnit_7.tgate_1.IN distortionUnit_7.myOpamp_0.INn VGND.t28 sky130_fd_pr__res_xhigh_po_0p69 l=10
X73 distortionUnit_3.tgate_1.IN distortionUnit_3.myOpamp_0.INn a_8014_30557# VGND.t276 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X74 bufferUnit_0.OUT ui_in[0].t2 bufferUnit_0.tgate_1.IN VGND.t174 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X75 a_20842_23723# distortionUnit_6.IN a_20584_23723# VGND.t273 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X76 a_8014_30557# a_6912_30102# VGND.t467 VGND.t379 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X77 VGND.t364 VGND.t362 VGND.t364 VGND.t363 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X78 distortionUnit_5.tgate_1.IN distortionUnit_5.myOpamp_0.INn a_8134_23853# VGND.t94 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X79 a_20842_23723# distortionUnit_6.IN a_20584_23723# VGND.t186 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X80 VGND.t361 VGND.t360 VGND.t361 VGND.t36 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X81 VGND.t359 VGND.t357 VGND.t359 VGND.t358 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X82 VGND.t10 ui_in[4].t4 distortionUnit_5.tgate_1.CTRLB VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X83 distortionUnit_2.tgate_1.IN distortionUnit_2.myOpamp_0.INn VGND.t39 sky130_fd_pr__res_xhigh_po_0p69 l=10
X84 distortionUnit_6.tgate_1.CTRLB ui_in[5].t2 VGND.t142 VGND.t141 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X85 distortionUnit_5.tgate_1.IN distortionUnit_5.myOpamp_0.INn a_8134_23853# VGND.t93 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X86 distortionUnit_3.IN ui_in[1].t3 bufferUnit_0.OUT VPWR.t46 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X87 bufferUnit_0.tgate_1.CTRLB ui_in[0].t3 VGND.t176 VGND.t175 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X88 a_7756_30557# VGND.t355 VGND.t356 VGND.t267 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X89 distortionUnit_6.tgate_1.IN distortionUnit_6.tgate_1.CTRLB distortionUnit_6.OUT VPWR.t56 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X90 VGND.t354 VGND.t352 VGND.t353 VGND.t323 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0 ps=0 w=0.42 l=1
X91 bufferUnit_0.tgate_1.CTRLB ui_in[0].t4 VGND.t178 VGND.t177 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X92 distortionUnit_4.tgate_1.IN ui_in[3].t4 distortionUnit_5.IN.t7 VGND.t163 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X93 a_20488_30481# distortionUnit_4.IN a_20746_30481# VGND.t43 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X94 VPWR.t178 a_20934_16677# a_20934_16677# VPWR.t177 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X95 distortionUnit_7.tgate_1.CTRLB ui_in[7].t1 VPWR.t91 distortionUnit_7.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X96 VPWR.t154 a_20488_30481# a_20488_30481# VPWR.t153 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X97 VGND.t351 VGND.t350 VGND.t351 VGND.t282 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X98 a_7756_30557# a_7756_30557# VPWR.t309 VPWR.t308 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X99 VPWR.t203 a_20584_23723# a_20584_23723# VPWR.t202 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X100 a_20584_23723# distortionUnit_6.IN a_20842_23723# VGND.t184 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X101 distortionUnit_4.tgate_1.IN distortionUnit_4.myOpamp_0.INn VGND.t153 sky130_fd_pr__res_xhigh_po_0p69 l=10
X102 bufferUnit_0.OUT bufferUnit_0.tgate_1.CTRLB bufferUnit_0.tgate_1.IN VPWR.t78 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X103 a_20934_16677# distortionUnit_7.IN a_21192_16677# VGND.t205 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X104 a_20584_23723# VGND.t348 VGND.t349 VGND.t257 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X105 distortionUnit_2.tgate_1.CTRLB ui_in[1].t4 VPWR.t47 distortionUnit_2.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X106 distortionUnit_4.tgate_1.CTRLB ui_in[3].t5 VGND.t165 VGND.t164 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X107 distortionUnit_0.tgate_1.IN a_7752_16807# VPWR.t128 VPWR.t127 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X108 VGND.t144 ui_in[5].t3 distortionUnit_6.tgate_1.CTRLB VGND.t143 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X109 VPWR.t43 ui_in[6].t5 distortionUnit_0.tgate_1.CTRLB distortionUnit_0.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X110 distortionUnit_7.tgate_1.CTRLB ui_in[7].t2 VPWR.t92 distortionUnit_7.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X111 VGND.t121 ui_in[0].t5 bufferUnit_0.tgate_1.CTRLB VGND.t120 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X112 VPWR.t93 ui_in[7].t3 distortionUnit_7.tgate_1.CTRLB distortionUnit_7.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X113 distortionUnit_0.tgate_1.IN distortionUnit_0.tgate_1.CTRLB distortionUnit_7.IN VPWR.t164 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X114 VGND.t347 VGND.t345 VGND.t347 VGND.t346 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X115 VGND.t344 VGND.t343 VGND.t344 VGND.t198 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X116 a_20746_30481# distortionUnit_4.myOpamp_0.INn distortionUnit_4.tgate_1.IN VGND.t154 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X117 distortionUnit_2.tgate_1.IN distortionUnit_2.myOpamp_0.INn a_20782_36601# VGND.t377 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X118 VPWR.t307 a_7756_30557# distortionUnit_3.tgate_1.IN VPWR.t306 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X119 VGND.t397 a_20090_16222# a_20090_16222# VGND.t197 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X120 a_7736_36483# a_7736_36483# VPWR.t227 VPWR.t226 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X121 VPWR.t44 ui_in[6].t6 distortionUnit_0.tgate_1.CTRLB distortionUnit_0.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X122 distortionUnit_3.tgate_1.CTRLB ui_in[2].t3 VPWR.t102 distortionUnit_3.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X123 a_8014_30557# distortionUnit_3.myOpamp_0.INn distortionUnit_3.tgate_1.IN VGND.t381 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X124 distortionUnit_2.tgate_1.CTRLB ui_in[1].t5 VPWR.t48 distortionUnit_2.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X125 bufferUnit_0.tgate_1.IN bufferUnit_0.tgate_1.IN a_7994_36483# VGND.t411 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X126 distortionUnit_2.tgate_1.IN a_20524_36601# VPWR.t74 VPWR.t73 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X127 VGND.t167 ui_in[3].t6 distortionUnit_4.tgate_1.CTRLB VGND.t166 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X128 VPWR.t108 a_19644_30026# VGND.t195 sky130_fd_pr__res_xhigh_po_0p35 l=0.16
X129 distortionUnit_6.OUT ui_in[5].t4 distortionUnit_6.tgate_1.IN VGND.t52 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X130 distortionUnit_2.tgate_1.IN a_20524_36601# VPWR.t70 VPWR.t69 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X131 a_20488_30481# a_20488_30481# VPWR.t152 VPWR.t151 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X132 a_20090_16222# a_20090_16222# VGND.t396 VGND.t202 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X133 a_19644_30026# a_19644_30026# VGND.t161 VGND.t40 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X134 a_20524_36601# bufferUnit_0.OUT a_20782_36601# VGND.t446 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X135 distortionUnit_3.tgate_1.CTRLB ui_in[2].t4 VPWR.t80 distortionUnit_3.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X136 VPWR.t81 ui_in[2].t5 distortionUnit_3.tgate_1.CTRLB distortionUnit_3.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X137 VGND.t342 VGND.t341 distortionUnit_6.tgate_1.IN VGND.t245 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X138 VGND.t340 VGND.t339 distortionUnit_5.tgate_1.IN VGND.t242 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X139 distortionUnit_7.tgate_1.IN distortionUnit_7.tgate_1.CTRLB ua[1].t5 VPWR.t286 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X140 VGND.t169 ui_in[3].t7 distortionUnit_4.tgate_1.CTRLB VGND.t168 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X141 distortionUnit_3.tgate_1.IN distortionUnit_3.myOpamp_0.INn a_8014_30557# VGND.t380 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X142 VPWR.t225 a_7736_36483# bufferUnit_0.tgate_1.IN VPWR.t224 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X143 bufferUnit_0.tgate_1.IN ui_in[0].t6 bufferUnit_0.OUT VGND.t122 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X144 a_20842_23723# distortionUnit_6.myOpamp_0.INn distortionUnit_6.tgate_1.IN VGND.t182 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X145 VPWR.t28 a_7876_23853# a_7876_23853# VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X146 distortionUnit_0.tgate_1.CTRLB ui_in[6].t7 VPWR.t45 distortionUnit_0.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X147 VGND.t338 VGND.t337 VGND.t338 VGND.t74 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X148 distortionUnit_3.tgate_1.IN distortionUnit_3.myOpamp_0.INn VGND.t179 sky130_fd_pr__res_xhigh_po_0p69 l=10
X149 distortionUnit_6.tgate_1.CTRLB ui_in[5].t5 VGND.t54 VGND.t53 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X150 VPWR.t176 a_20934_16677# a_20934_16677# VPWR.t175 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X151 distortionUnit_3.tgate_1.IN distortionUnit_3.myOpamp_0.INn a_8014_30557# VGND.t239 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X152 VGND.t106 a_6908_16352# a_6908_16352# VGND.t105 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X153 VPWR.t72 a_20524_36601# a_20524_36601# VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X154 a_8134_23853# distortionUnit_5.IN.t12 a_7876_23853# VGND.t236 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X155 distortionUnit_7.IN ui_in[6].t8 distortionUnit_0.tgate_1.IN VGND.t65 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X156 VPWR.t68 a_20524_36601# a_20524_36601# VPWR.t67 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X157 bufferUnit_0.tgate_1.CTRLB ui_in[0].t7 VGND.t124 VGND.t123 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X158 distortionUnit_0.tgate_1.IN distortionUnit_0.myOpamp_0.INn VGND.t23 sky130_fd_pr__res_xhigh_po_0p69 l=10
X159 VPWR.t150 a_20488_30481# distortionUnit_4.tgate_1.IN VPWR.t149 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X160 a_20782_36601# distortionUnit_2.myOpamp_0.INn distortionUnit_2.tgate_1.IN VGND.t407 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X161 VGND.t336 VGND.t334 VGND.t335 VGND.t248 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0 ps=0 w=0.42 l=1
X162 distortionUnit_4.tgate_1.IN distortionUnit_4.tgate_1.CTRLB distortionUnit_5.IN.t11 VPWR.t207 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X163 ua[1].t4 distortionUnit_7.tgate_1.CTRLB distortionUnit_7.tgate_1.IN VPWR.t285 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X164 VGND.t333 VGND.t331 distortionUnit_0.tgate_1.IN VGND.t332 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X165 VGND.t136 ui_in[2].t6 distortionUnit_3.tgate_1.CTRLB VGND.t135 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X166 VGND.t330 VGND.t328 VGND.t330 VGND.t329 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X167 a_8010_16807# distortionUnit_6.OUT a_7752_16807# VGND.t107 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X168 a_20934_16677# VPWR.t262 VPWR.t264 VPWR.t263 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X169 distortionUnit_6.tgate_1.CTRLB ui_in[5].t6 VGND.t56 VGND.t55 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X170 VGND.t466 a_6912_30102# a_8014_30557# VGND.t73 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X171 VPWR.t51 a_7032_23398# VGND.t72 sky130_fd_pr__res_xhigh_po_0p35 l=0.16
X172 VGND.t327 VGND.t325 VGND.t327 VGND.t326 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X173 bufferUnit_0.tgate_1.CTRLB ui_in[0].t8 VGND.t126 VGND.t125 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X174 VGND.t58 ui_in[5].t7 distortionUnit_6.tgate_1.CTRLB VGND.t57 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X175 VGND.t69 ui_in[0].t9 bufferUnit_0.tgate_1.CTRLB VGND.t68 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X176 distortionUnit_7.tgate_1.CTRLB ui_in[7].t4 VPWR.t94 distortionUnit_7.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X177 a_20524_36601# VPWR.t259 VPWR.t261 VPWR.t260 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X178 VPWR.t82 ui_in[7].t5 distortionUnit_7.tgate_1.CTRLB distortionUnit_7.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X179 VPWR.t107 a_19680_36146# VGND.t194 sky130_fd_pr__res_xhigh_po_0p35 l=0.16
X180 distortionUnit_7.IN distortionUnit_0.tgate_1.CTRLB distortionUnit_0.tgate_1.IN VPWR.t163 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X181 distortionUnit_0.tgate_1.IN distortionUnit_0.myOpamp_0.INn a_8010_16807# VGND.t358 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X182 distortionUnit_5.IN.t9 distortionUnit_4.tgate_1.CTRLB distortionUnit_4.IN VGND.t421 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X183 distortionUnit_3.tgate_1.CTRLB ui_in[2].t7 VGND.t138 VGND.t137 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X184 VPWR.t126 a_7752_16807# a_7752_16807# VPWR.t125 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X185 VPWR.t83 ui_in[7].t6 distortionUnit_7.tgate_1.CTRLB distortionUnit_7.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X186 distortionUnit_6.tgate_1.IN distortionUnit_6.myOpamp_0.INn VGND.t438 sky130_fd_pr__res_xhigh_po_0p69 l=10
X187 VGND.t191 a_19740_23268# a_20842_23723# VGND.t190 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X188 VPWR.t96 ui_in[3].t8 distortionUnit_4.tgate_1.CTRLB distortionUnit_4.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X189 distortionUnit_4.tgate_1.IN distortionUnit_4.myOpamp_0.INn a_20746_30481# VGND.t227 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X190 ua[1].t1 ui_in[7].t7 distortionUnit_7.tgate_1.IN VGND.t139 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X191 a_21192_16677# distortionUnit_7.IN a_20934_16677# VGND.t204 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X192 distortionUnit_3.tgate_1.CTRLB ui_in[2].t8 VGND.t25 VGND.t24 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X193 VGND.t417 a_6892_36028# a_7994_36483# VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X194 distortionUnit_5.tgate_1.IN distortionUnit_5.myOpamp_0.INn VGND.t192 sky130_fd_pr__res_xhigh_po_0p69 l=10
X195 VPWR.t305 a_7756_30557# a_7756_30557# VPWR.t304 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X196 a_7752_16807# VGND.t322 VGND.t324 VGND.t323 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X197 VGND.t314 VGND.t313 bufferUnit_0.tgate_1.IN VGND.t222 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X198 distortionUnit_2.tgate_1.CTRLB ui_in[1].t6 VPWR.t109 distortionUnit_2.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X199 distortionUnit_0.tgate_1.CTRLB ui_in[6].t9 VGND.t67 VGND.t66 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X200 VGND.t321 VGND.t320 VGND.t321 VGND.t201 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X201 VPWR.t110 ui_in[1].t7 distortionUnit_2.tgate_1.CTRLB distortionUnit_2.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X202 a_7876_23853# distortionUnit_5.IN.t13 a_8134_23853# VGND.t146 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X203 VGND.t444 a_19680_36146# a_20782_36601# VGND.t443 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X204 VGND.t319 VGND.t318 VGND.t319 VGND.t233 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X205 a_7994_36483# ua[0].t6 a_7736_36483# VGND.t409 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X206 VPWR.t84 ui_in[7].t8 distortionUnit_7.tgate_1.CTRLB distortionUnit_7.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X207 distortionUnit_7.tgate_1.CTRLB ui_in[7].t9 VPWR.t85 distortionUnit_7.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X208 a_20746_30481# a_19644_30026# VGND.t160 VGND.t159 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X209 a_7994_36483# ua[0].t7 a_7736_36483# VGND.t219 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X210 distortionUnit_2.tgate_1.IN distortionUnit_2.tgate_1.CTRLB distortionUnit_3.IN VPWR.t98 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X211 VPWR.t124 a_7752_16807# distortionUnit_0.tgate_1.IN VPWR.t123 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X212 distortionUnit_7.tgate_1.IN ui_in[7].t10 ua[1].t0 VGND.t109 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X213 a_20842_23723# a_19740_23268# VGND.t189 VGND.t188 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X214 VPWR.t9 ui_in[4].t5 distortionUnit_5.tgate_1.CTRLB distortionUnit_5.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X215 VPWR.t111 ui_in[1].t8 distortionUnit_2.tgate_1.CTRLB distortionUnit_2.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X216 VPWR.t174 a_20934_16677# distortionUnit_7.tgate_1.IN VPWR.t173 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X217 distortionUnit_4.tgate_1.CTRLB ui_in[3].t9 VPWR.t157 distortionUnit_4.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X218 bufferUnit_0.tgate_1.IN bufferUnit_0.tgate_1.IN a_7994_36483# VGND.t213 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X219 a_7994_36483# a_6892_36028# VGND.t416 VGND.t415 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X220 VGND.t317 VGND.t315 VGND.t316 VGND.t230 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0 ps=0 w=0.42 l=1
X221 VPWR.t33 ui_in[2].t9 distortionUnit_3.tgate_1.CTRLB distortionUnit_3.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X222 a_7756_30557# a_7756_30557# VPWR.t303 VPWR.t302 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X223 distortionUnit_6.tgate_1.IN distortionUnit_6.myOpamp_0.INn a_20842_23723# VGND.t180 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X224 VPWR.t66 a_20524_36601# distortionUnit_2.tgate_1.IN VPWR.t65 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X225 VPWR.t10 ui_in[1].t9 distortionUnit_2.tgate_1.CTRLB distortionUnit_2.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X226 VPWR.t223 a_7736_36483# a_7736_36483# VPWR.t222 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X227 a_8134_23853# distortionUnit_5.myOpamp_0.INn distortionUnit_5.tgate_1.IN VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X228 a_8014_30557# distortionUnit_3.IN a_7756_30557# VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X229 VPWR.t106 a_6892_36028# VGND.t193 sky130_fd_pr__res_xhigh_po_0p35 l=0.16
X230 distortionUnit_3.IN distortionUnit_2.tgate_1.CTRLB bufferUnit_0.OUT VGND.t171 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X231 distortionUnit_3.IN distortionUnit_2.tgate_1.CTRLB distortionUnit_2.tgate_1.IN VPWR.t97 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X232 a_7736_36483# VGND.t311 VGND.t312 VGND.t207 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X233 distortionUnit_0.tgate_1.IN ui_in[6].t10 distortionUnit_7.IN VGND.t427 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X234 distortionUnit_7.tgate_1.CTRLB ui_in[7].t11 VGND.t111 VGND.t110 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X235 distortionUnit_0.tgate_1.IN a_7752_16807# VPWR.t122 VPWR.t121 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X236 VPWR.t162 a_20090_16222# VGND.t382 sky130_fd_pr__res_xhigh_po_0p35 l=0.16
X237 VGND.t310 VGND.t308 VGND.t310 VGND.t309 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X238 a_20746_30481# distortionUnit_4.IN a_20488_30481# VGND.t42 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X239 VPWR.t34 ui_in[2].t10 distortionUnit_3.tgate_1.CTRLB distortionUnit_3.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X240 VPWR a_6908_16352# VGND sky130_fd_pr__res_xhigh_po_0p35 l=26.11
X241 distortionUnit_4.tgate_1.IN a_20488_30481# VPWR.t148 VPWR.t147 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X242 distortionUnit_6.tgate_1.IN a_20584_23723# VPWR.t201 VPWR.t200 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X243 distortionUnit_5.IN.t4 ui_in[3].t10 distortionUnit_4.IN VPWR.t158 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X244 VGND distortionUnit_0.myOpamp_0.INn VGND.t383 sky130_fd_pr__res_xhigh_po_0p69 l=4
X245 distortionUnit_7.tgate_1.IN a_20934_16677# VPWR.t172 VPWR.t171 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X246 VGND.t307 VGND.t306 VGND.t307 VGND.t261 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X247 VPWR.t95 a_6912_30102# VGND.t152 sky130_fd_pr__res_xhigh_po_0p35 l=0.16
X248 VGND.t401 ui_in[5].t8 distortionUnit_6.tgate_1.CTRLB VGND.t400 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X249 a_20842_23723# distortionUnit_6.IN a_20584_23723# VGND.t370 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X250 a_7032_23398# a_7032_23398# VGND.t151 VGND.t37 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X251 distortionUnit_7.tgate_1.CTRLB ui_in[7].t12 VGND.t113 VGND.t112 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X252 a_7736_36483# a_7736_36483# VPWR.t221 VPWR.t220 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X253 bufferUnit_0.OUT distortionUnit_2.tgate_1.CTRLB distortionUnit_3.IN VGND.t170 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X254 VGND.t115 ui_in[7].t13 distortionUnit_7.tgate_1.CTRLB VGND.t114 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X255 a_8010_16807# a_6908_16352# VGND.t104 VGND.t103 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X256 VGND.t71 ui_in[0].t10 bufferUnit_0.tgate_1.CTRLB VGND.t70 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X257 a_20584_23723# a_20584_23723# VPWR.t199 VPWR.t198 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X258 distortionUnit_0.tgate_1.IN distortionUnit_0.myOpamp_0.INn a_8010_16807# VGND.t105 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X259 a_20488_30481# distortionUnit_4.IN a_20746_30481# VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X260 a_21192_16677# a_20090_16222# VGND.t395 VGND.t196 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X261 VGND.t403 ui_in[5].t9 distortionUnit_6.tgate_1.CTRLB VGND.t402 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X262 VGND.t305 VGND.t304 VGND.t305 VGND.t91 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X263 distortionUnit_3.tgate_1.CTRLB ui_in[2].t11 VGND.t27 VGND.t26 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X264 distortionUnit_0.tgate_1.CTRLB ui_in[6].t11 VGND.t429 VGND.t428 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X265 VGND.t150 a_7032_23398# a_8134_23853# VGND.t38 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X266 a_7756_30557# distortionUnit_3.IN a_8014_30557# VGND.t75 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X267 VGND distortionUnit_6.myOpamp_0.INn VGND.t469 sky130_fd_pr__res_xhigh_po_0p69 l=4
X268 a_7994_36483# bufferUnit_0.tgate_1.IN bufferUnit_0.tgate_1.IN VGND.t418 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X269 a_20934_16677# distortionUnit_7.IN a_21192_16677# VGND.t203 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X270 VGND.t303 VGND.t300 VGND.t302 VGND.t301 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0 ps=0 w=0.42 l=1
X271 VGND distortionUnit_4.myOpamp_0.INn VGND.t62 sky130_fd_pr__res_xhigh_po_0p69 l=4
X272 VPWR a_19740_23268# VGND sky130_fd_pr__res_xhigh_po_0p35 l=26.11
X273 distortionUnit_3.tgate_1.CTRLB ui_in[2].t12 VGND.t81 VGND.t80 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X274 VGND.t299 VGND.t297 VGND.t299 VGND.t298 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X275 VPWR.t146 a_20488_30481# a_20488_30481# VPWR.t145 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X276 VGND.t83 ui_in[2].t13 distortionUnit_3.tgate_1.CTRLB VGND.t82 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X277 VGND.t158 a_19644_30026# a_19644_30026# VGND.t157 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X278 a_20782_36601# bufferUnit_0.OUT a_20524_36601# VGND.t326 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X279 VPWR.t159 ui_in[3].t11 distortionUnit_4.tgate_1.CTRLB distortionUnit_4.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X280 VPWR.t197 a_20584_23723# distortionUnit_6.tgate_1.IN VPWR.t196 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X281 distortionUnit_6.IN ui_in[4].t6 distortionUnit_5.IN.t1 VPWR.t8 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X282 VGND.t431 ui_in[6].t12 distortionUnit_0.tgate_1.CTRLB VGND.t430 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X283 distortionUnit_4.tgate_1.CTRLB ui_in[3].t12 VPWR.t160 distortionUnit_4.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X284 VGND.t296 VGND.t295 VGND.t296 VGND.t200 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X285 distortionUnit_6.tgate_1.CTRLB ui_in[5].t10 VGND.t405 VGND.t404 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X286 a_21192_16677# distortionUnit_7.myOpamp_0.INn distortionUnit_7.tgate_1.IN VGND.t199 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X287 VGND.t433 ui_in[6].t13 distortionUnit_0.tgate_1.CTRLB VGND.t432 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X288 VPWR.t11 ui_in[1].t10 distortionUnit_2.tgate_1.CTRLB distortionUnit_2.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X289 VGND.t294 VGND.t292 VGND.t294 VGND.t293 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X290 a_8014_30557# distortionUnit_3.myOpamp_0.INn distortionUnit_3.tgate_1.IN VGND.t379 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X291 distortionUnit_2.tgate_1.CTRLB ui_in[1].t11 VPWR.t12 distortionUnit_2.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X292 bufferUnit_0.tgate_1.IN bufferUnit_0.tgate_1.IN a_7994_36483# VGND.t363 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X293 a_8134_23853# distortionUnit_5.IN.t14 a_7876_23853# VGND.t36 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X294 distortionUnit_2.tgate_1.IN a_20524_36601# VPWR.t64 VPWR.t63 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X295 a_20488_30481# a_20488_30481# VPWR.t144 VPWR.t143 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X296 distortionUnit_5.IN.t3 distortionUnit_5.tgate_1.CTRLB distortionUnit_6.IN VGND.t79 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X297 distortionUnit_6.tgate_1.CTRLB ui_in[5].t11 VPWR.t185 distortionUnit_6.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X298 VGND.t291 VGND.t290 VGND.t291 VGND.t44 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X299 a_20524_36601# bufferUnit_0.OUT a_20782_36601# VGND.t443 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X300 distortionUnit_4.tgate_1.CTRLB ui_in[3].t13 VPWR.t161 distortionUnit_4.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X301 distortionUnit_0.tgate_1.CTRLB ui_in[6].t14 VGND.t435 VGND.t434 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X302 distortionUnit_5.tgate_1.CTRLB ui_in[4].t7 VPWR.t7 distortionUnit_5.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X303 VGND.t289 VGND.t287 VGND.t289 VGND.t288 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X304 VGND.t286 VGND.t284 VGND.t286 VGND.t285 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X305 VPWR.t49 ui_in[0].t11 bufferUnit_0.tgate_1.CTRLB bufferUnit_0.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X306 VGND.t283 VGND.t281 distortionUnit_7.tgate_1.IN VGND.t282 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X307 a_20934_16677# a_20934_16677# VPWR.t170 VPWR.t169 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X308 a_8134_23853# a_7032_23398# VGND.t149 VGND.t95 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X309 VPWR.t26 a_7876_23853# a_7876_23853# VPWR.t25 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X310 distortionUnit_7.tgate_1.CTRLB ui_in[7].t14 VGND.t117 VGND.t116 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X311 a_6912_30102# a_6912_30102# VGND.t465 VGND.t77 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X312 bufferUnit_0.tgate_1.IN a_7736_36483# VPWR.t219 VPWR.t218 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X313 VGND.t280 VGND.t278 VGND.t280 VGND.t279 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X314 VGND.t414 a_6892_36028# a_7994_36483# VGND.t413 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X315 VGND.t128 ui_in[7].t15 distortionUnit_7.tgate_1.CTRLB VGND.t127 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X316 a_20524_36601# a_20524_36601# VPWR.t62 VPWR.t61 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X317 VGND.t442 a_19680_36146# a_19680_36146# VGND.t406 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X318 distortionUnit_5.tgate_1.CTRLB ui_in[4].t8 VPWR.t6 distortionUnit_5.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X319 VGND.t130 ui_in[7].t16 distortionUnit_7.tgate_1.CTRLB VGND.t129 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X320 VGND distortionUnit_3.myOpamp_0.INn VGND.t59 sky130_fd_pr__res_xhigh_po_0p69 l=4
X321 VPWR a_6892_36028# VGND sky130_fd_pr__res_xhigh_po_0p35 l=26.11
X322 VPWR.t5 ui_in[4].t9 distortionUnit_5.tgate_1.CTRLB distortionUnit_5.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X323 VPWR.t120 a_7752_16807# a_7752_16807# VPWR.t119 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X324 distortionUnit_5.tgate_1.IN a_7876_23853# VPWR.t24 VPWR.t23 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X325 VPWR.t288 ui_in[5].t12 distortionUnit_6.tgate_1.CTRLB distortionUnit_6.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X326 VGND.t277 VGND.t275 VGND.t277 VGND.t276 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X327 bufferUnit_0.tgate_1.CTRLB ui_in[0].t12 VPWR.t50 bufferUnit_0.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X328 VGND.t274 VGND.t272 VGND.t274 VGND.t273 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X329 distortionUnit_7.tgate_1.IN distortionUnit_7.myOpamp_0.INn a_21192_16677# VGND.t198 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X330 distortionUnit_4.tgate_1.IN distortionUnit_4.myOpamp_0.INn a_20746_30481# VGND.t346 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X331 distortionUnit_3.IN ui_in[2].t14 distortionUnit_4.IN VPWR.t54 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X332 VGND.t148 a_7032_23398# a_7032_23398# VGND.t94 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X333 a_7876_23853# a_7876_23853# VPWR.t22 VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X334 distortionUnit_6.OUT ui_in[5].t13 distortionUnit_6.IN VPWR.t289 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X335 a_19740_23268# a_19740_23268# VGND.t187 VGND.t186 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X336 distortionUnit_6.IN distortionUnit_5.tgate_1.CTRLB distortionUnit_5.tgate_1.IN VPWR.t53 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X337 a_8010_16807# distortionUnit_6.OUT a_7752_16807# VGND.t309 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X338 bufferUnit_0.tgate_1.CTRLB ui_in[0].t13 VPWR.t86 bufferUnit_0.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X339 distortionUnit_7.tgate_1.IN distortionUnit_7.myOpamp_0.INn a_21192_16677# VGND.t197 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X340 VGND.t271 VGND.t270 VGND.t271 VGND.t93 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X341 a_7876_23853# VPWR.t256 VPWR.t258 VPWR.t257 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X342 VGND.t132 ui_in[7].t17 distortionUnit_7.tgate_1.CTRLB VGND.t131 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X343 VGND.t269 VGND.t266 VGND.t268 VGND.t267 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0 ps=0 w=0.42 l=1
X344 a_19680_36146# a_19680_36146# VGND.t441 VGND.t440 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X345 distortionUnit_7.tgate_1.CTRLB ui_in[7].t18 VGND.t134 VGND.t133 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X346 VPWR.t60 a_20524_36601# distortionUnit_2.tgate_1.IN VPWR.t59 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X347 VGND.t265 VGND.t263 VGND.t265 VGND.t264 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X348 VGND.t262 VGND.t260 distortionUnit_2.tgate_1.IN VGND.t261 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X349 a_7752_16807# a_7752_16807# VPWR.t118 VPWR.t117 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X350 VPWR.t4 ui_in[4].t10 distortionUnit_5.tgate_1.CTRLB distortionUnit_5.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X351 VGND.t156 a_19644_30026# a_20746_30481# VGND.t43 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X352 distortionUnit_5.IN.t6 ui_in[3].t14 distortionUnit_4.tgate_1.IN VGND.t33 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X353 VGND.t8 ui_in[4].t11 distortionUnit_5.tgate_1.CTRLB VGND.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X354 distortionUnit_4.tgate_1.CTRLB ui_in[3].t15 VPWR.t36 distortionUnit_4.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X355 a_7752_16807# a_7752_16807# VPWR.t116 VPWR.t115 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X356 distortionUnit_4.IN distortionUnit_3.tgate_1.CTRLB distortionUnit_3.IN VGND.t456 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X357 VPWR.t255 VPWR.t253 distortionUnit_3.tgate_1.IN VPWR.t254 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X358 distortionUnit_6.IN distortionUnit_6.tgate_1.CTRLB distortionUnit_6.OUT VGND.t87 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X359 VPWR.t41 a_6908_16352# VGND.t51 sky130_fd_pr__res_xhigh_po_0p35 l=0.16
X360 VPWR.t87 ui_in[0].t14 bufferUnit_0.tgate_1.CTRLB bufferUnit_0.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X361 VGND.t185 a_19740_23268# a_20842_23723# VGND.t184 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X362 VGND.t85 ui_in[2].t15 distortionUnit_3.tgate_1.CTRLB VGND.t84 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X363 distortionUnit_5.tgate_1.IN ui_in[4].t12 distortionUnit_6.IN VGND.t6 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X364 distortionUnit_2.tgate_1.CTRLB ui_in[1].t12 VGND.t423 VGND.t422 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X365 a_21192_16677# distortionUnit_7.IN a_20934_16677# VGND.t202 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X366 a_8010_16807# distortionUnit_0.myOpamp_0.INn distortionUnit_0.tgate_1.IN VGND.t103 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X367 a_20746_30481# distortionUnit_4.IN a_20488_30481# VGND.t40 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X368 VPWR.t301 a_7756_30557# a_7756_30557# VPWR.t300 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X369 VGND.t394 a_20090_16222# a_21192_16677# VGND.t205 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X370 VGND.t437 ui_in[6].t15 distortionUnit_0.tgate_1.CTRLB VGND.t436 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X371 VGND.t259 VGND.t256 VGND.t258 VGND.t257 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0 ps=0 w=0.42 l=1
X372 distortionUnit_3.tgate_1.IN distortionUnit_3.tgate_1.CTRLB distortionUnit_4.IN VPWR.t280 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X373 ua[0].t3 ui_in[0].t15 bufferUnit_0.OUT VPWR.t88 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X374 VGND distortionUnit_7.myOpamp_0.INn VGND.t389 sky130_fd_pr__res_xhigh_po_0p69 l=4
X375 VGND.t255 VGND.t253 VGND.t254 VGND.t216 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0 ps=0 w=0.42 l=1
X376 a_8014_30557# distortionUnit_3.IN a_7756_30557# VGND.t74 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X377 VGND.t30 ui_in[2].t16 distortionUnit_3.tgate_1.CTRLB VGND.t29 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X378 a_20746_30481# a_19644_30026# VGND.t155 VGND.t154 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X379 VPWR.t114 a_7752_16807# distortionUnit_0.tgate_1.IN VPWR.t113 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X380 VPWR a_19644_30026# VGND sky130_fd_pr__res_xhigh_po_0p35 l=26.11
X381 VGND.t252 VGND.t250 VGND.t252 VGND.t251 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X382 distortionUnit_6.tgate_1.CTRLB ui_in[5].t14 VPWR.t290 distortionUnit_6.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X383 distortionUnit_3.tgate_1.IN a_7756_30557# VPWR.t299 VPWR.t298 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X384 VGND.t48 ui_in[6].t16 distortionUnit_0.tgate_1.CTRLB VGND.t47 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X385 distortionUnit_4.tgate_1.IN a_20488_30481# VPWR.t142 VPWR.t141 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X386 VPWR.t37 ui_in[3].t16 distortionUnit_4.tgate_1.CTRLB distortionUnit_4.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X387 distortionUnit_6.tgate_1.IN a_20584_23723# VPWR.t195 VPWR.t194 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X388 distortionUnit_5.IN.t10 distortionUnit_4.tgate_1.CTRLB distortionUnit_4.tgate_1.IN VPWR.t206 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X389 distortionUnit_2.tgate_1.CTRLB ui_in[1].t13 VGND.t425 VGND.t424 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X390 VPWR.t20 a_7876_23853# distortionUnit_5.tgate_1.IN VPWR.t19 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X391 distortionUnit_0.tgate_1.IN distortionUnit_0.myOpamp_0.INn a_8010_16807# VGND.t298 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X392 a_20488_30481# VGND.t247 VGND.t249 VGND.t248 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X393 VPWR.t252 VPWR.t250 bufferUnit_0.tgate_1.IN VPWR.t251 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X394 bufferUnit_0.OUT bufferUnit_0.tgate_1.CTRLB ua[0].t1 VGND.t119 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X395 a_8014_30557# a_6912_30102# VGND.t464 VGND.t381 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X396 a_7756_30557# VPWR.t247 VPWR.t249 VPWR.t248 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X397 VGND.t412 a_6892_36028# a_6892_36028# VGND.t411 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X398 distortionUnit_6.tgate_1.IN distortionUnit_6.myOpamp_0.INn a_20842_23723# VGND.t329 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X399 VPWR a_7032_23398# VGND sky130_fd_pr__res_xhigh_po_0p35 l=26.11
X400 VPWR.t217 a_7736_36483# a_7736_36483# VPWR.t216 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X401 distortionUnit_5.tgate_1.CTRLB ui_in[4].t13 VPWR.t3 distortionUnit_5.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X402 a_7756_30557# distortionUnit_3.IN a_8014_30557# VGND.t73 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X403 VPWR.t215 a_7736_36483# a_7736_36483# VPWR.t214 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X404 distortionUnit_3.IN ui_in[1].t14 distortionUnit_2.tgate_1.IN VGND.t426 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X405 VPWR.t38 ui_in[3].t17 distortionUnit_4.tgate_1.CTRLB distortionUnit_4.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X406 VGND.t102 a_6908_16352# a_8010_16807# VGND.t101 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X407 distortionUnit_6.tgate_1.CTRLB ui_in[5].t15 VPWR.t291 distortionUnit_6.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X408 VGND.t246 VGND.t244 VGND.t246 VGND.t245 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X409 VPWR.t193 a_20584_23723# a_20584_23723# VPWR.t192 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X410 VGND.t100 a_6908_16352# a_8010_16807# VGND.t99 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X411 VPWR.t133 ui_in[5].t16 distortionUnit_6.tgate_1.CTRLB distortionUnit_6.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X412 distortionUnit_4.IN distortionUnit_4.tgate_1.CTRLB distortionUnit_5.IN.t8 VGND.t420 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X413 distortionUnit_0.tgate_1.CTRLB ui_in[6].t17 VGND.t50 VGND.t49 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X414 distortionUnit_5.tgate_1.CTRLB ui_in[4].t14 VPWR.t2 distortionUnit_5.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X415 distortionUnit_5.tgate_1.IN a_7876_23853# VPWR.t18 VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X416 VPWR.t168 a_20934_16677# a_20934_16677# VPWR.t167 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X417 VGND.t243 VGND.t241 VGND.t243 VGND.t242 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X418 VPWR.t140 a_20488_30481# a_20488_30481# VPWR.t139 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X419 bufferUnit_0.tgate_1.IN a_7736_36483# VPWR.t213 VPWR.t212 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X420 VGND.t463 a_6912_30102# a_6912_30102# VGND.t380 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X421 a_20842_23723# a_19740_23268# VGND.t183 VGND.t182 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X422 VPWR.t191 a_20584_23723# a_20584_23723# VPWR.t190 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X423 distortionUnit_4.IN ui_in[2].t17 distortionUnit_3.IN VPWR.t35 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X424 bufferUnit_0.tgate_1.CTRLB ui_in[0].t16 VPWR.t89 bufferUnit_0.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X425 distortionUnit_5.tgate_1.IN a_7876_23853# VPWR.t16 VPWR.t15 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X426 distortionUnit_4.IN ui_in[2].t18 distortionUnit_3.tgate_1.IN VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X427 a_20584_23723# distortionUnit_6.IN a_20842_23723# VGND.t190 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X428 VGND.t240 VGND.t238 VGND.t240 VGND.t239 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X429 a_20782_36601# a_19680_36146# VGND.t439 VGND.t408 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X430 a_7736_36483# ua[0].t8 a_7994_36483# VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X431 VGND.t237 VGND.t235 VGND.t237 VGND.t236 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X432 distortionUnit_2.tgate_1.IN ui_in[1].t15 distortionUnit_3.IN VGND.t18 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X433 a_7736_36483# VPWR.t244 VPWR.t246 VPWR.t245 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X434 a_21192_16677# distortionUnit_7.IN a_20934_16677# VGND.t201 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X435 VPWR.t1 ui_in[4].t15 distortionUnit_5.tgate_1.CTRLB distortionUnit_5.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X436 VGND.t35 ui_in[3].t18 distortionUnit_4.tgate_1.CTRLB VGND.t34 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X437 a_8010_16807# a_6908_16352# VGND.t98 VGND.t97 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X438 distortionUnit_0.tgate_1.CTRLB ui_in[6].t18 VPWR.t39 distortionUnit_0.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X439 distortionUnit_6.IN ui_in[5].t17 distortionUnit_6.OUT VPWR.t134 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X440 VGND.t234 VGND.t232 distortionUnit_4.tgate_1.IN VGND.t233 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X441 distortionUnit_2.tgate_1.IN distortionUnit_2.myOpamp_0.INn a_20782_36601# VGND.t279 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X442 bufferUnit_0.tgate_1.CTRLB ui_in[0].t17 VPWR.t103 bufferUnit_0.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X443 a_20584_23723# a_20584_23723# VPWR.t189 VPWR.t188 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X444 VPWR.t104 ui_in[0].t18 bufferUnit_0.tgate_1.CTRLB bufferUnit_0.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X445 distortionUnit_5.IN.t0 ui_in[4].t16 distortionUnit_6.IN VPWR.t0 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X446 a_20746_30481# distortionUnit_4.myOpamp_0.INn distortionUnit_4.tgate_1.IN VGND.t159 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X447 distortionUnit_2.tgate_1.IN distortionUnit_2.myOpamp_0.INn a_20782_36601# VGND.t406 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X448 a_20488_30481# VPWR.t241 VPWR.t243 VPWR.t242 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X449 distortionUnit_3.IN distortionUnit_3.tgate_1.CTRLB distortionUnit_4.IN VGND.t455 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X450 VPWR.t297 a_7756_30557# distortionUnit_3.tgate_1.IN VPWR.t296 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X451 a_20584_23723# VPWR.t238 VPWR.t240 VPWR.t239 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X452 a_20842_23723# distortionUnit_6.myOpamp_0.INn distortionUnit_6.tgate_1.IN VGND.t188 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X453 distortionUnit_4.IN distortionUnit_3.tgate_1.CTRLB distortionUnit_3.tgate_1.IN VPWR.t279 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X454 bufferUnit_0.OUT ui_in[0].t19 ua[0].t2 VPWR.t105 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X455 a_7994_36483# bufferUnit_0.tgate_1.IN bufferUnit_0.tgate_1.IN VGND.t415 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X456 a_20934_16677# VGND.t229 VGND.t231 VGND.t230 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X457 distortionUnit_6.OUT distortionUnit_6.tgate_1.CTRLB distortionUnit_6.IN VGND.t86 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X458 distortionUnit_4.tgate_1.CTRLB ui_in[3].t19 VGND.t46 VGND.t45 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X459 distortionUnit_6.OUT ui_in[6].t19 distortionUnit_7.IN VPWR.t40 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X460 distortionUnit_5.tgate_1.CTRLB ui_in[4].t17 VGND.t5 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X461 distortionUnit_6.IN distortionUnit_5.tgate_1.CTRLB distortionUnit_5.IN.t2 VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X462 VGND.t228 VGND.t226 VGND.t228 VGND.t227 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X463 a_20782_36601# bufferUnit_0.OUT a_20524_36601# VGND.t440 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X464 distortionUnit_3.tgate_1.IN a_7756_30557# VPWR.t295 VPWR.t294 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X465 VGND.t225 VGND.t224 VGND.t225 VGND.t204 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X466 distortionUnit_2.tgate_1.CTRLB ui_in[1].t16 VGND.t20 VGND.t19 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X467 VGND.t22 ui_in[1].t17 distortionUnit_2.tgate_1.CTRLB VGND.t21 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X468 a_20782_36601# bufferUnit_0.OUT a_20524_36601# VGND.t264 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X469 VGND distortionUnit_2.myOpamp_0.INn VGND.t386 sky130_fd_pr__res_xhigh_po_0p69 l=4
X470 distortionUnit_3.tgate_1.IN a_7756_30557# VPWR.t293 VPWR.t292 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X471 VGND.t223 VGND.t221 VGND.t223 VGND.t222 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X472 VGND.t147 a_7032_23398# a_8134_23853# VGND.t146 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X473 VPWR.t211 a_7736_36483# bufferUnit_0.tgate_1.IN VPWR.t210 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X474 ua[0].t0 bufferUnit_0.tgate_1.CTRLB bufferUnit_0.OUT VGND.t118 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X475 a_6892_36028# a_6892_36028# VGND.t410 VGND.t409 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X476 distortionUnit_5.tgate_1.CTRLB ui_in[4].t18 VGND.t3 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X477 VPWR.t58 a_20524_36601# a_20524_36601# VPWR.t57 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X478 VGND.t1 ui_in[4].t19 distortionUnit_5.tgate_1.CTRLB VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X479 VGND.t220 VGND.t218 VGND.t220 VGND.t219 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X480 a_8134_23853# distortionUnit_5.IN.t15 a_7876_23853# VGND.t37 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X481 distortionUnit_7.IN distortionUnit_0.tgate_1.CTRLB distortionUnit_6.OUT VGND.t392 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X482 VPWR.t237 VPWR.t235 distortionUnit_4.tgate_1.IN VPWR.t236 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X483 VPWR.t234 VPWR.t232 distortionUnit_6.tgate_1.IN VPWR.t233 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X484 VGND.t473 ui_in[1].t18 distortionUnit_2.tgate_1.CTRLB VGND.t472 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X485 VPWR.t135 ui_in[5].t18 distortionUnit_6.tgate_1.CTRLB distortionUnit_6.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X486 VPWR.t231 VPWR.t229 distortionUnit_5.tgate_1.IN VPWR.t230 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X487 VPWR.t138 a_20488_30481# distortionUnit_4.tgate_1.IN VPWR.t137 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X488 a_20524_36601# VGND.t215 VGND.t217 VGND.t216 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X489 VPWR.t187 a_20584_23723# distortionUnit_6.tgate_1.IN VPWR.t186 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X490 VPWR a_20090_16222# VGND sky130_fd_pr__res_xhigh_po_0p35 l=26.11
X491 VGND.t214 VGND.t212 VGND.t214 VGND.t213 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X492 VGND.t475 ui_in[1].t19 distortionUnit_2.tgate_1.CTRLB VGND.t474 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X493 distortionUnit_6.OUT distortionUnit_6.tgate_1.CTRLB distortionUnit_6.tgate_1.IN VPWR.t55 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X494 distortionUnit_5.tgate_1.IN distortionUnit_5.tgate_1.CTRLB distortionUnit_6.IN VPWR.t52 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X495 distortionUnit_7.IN ui_in[7].t19 ua[1].t2 VPWR.t77 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X496 VGND.t181 a_19740_23268# a_19740_23268# VGND.t180 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X497 a_21192_16677# distortionUnit_7.myOpamp_0.INn distortionUnit_7.tgate_1.IN VGND.t196 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X498 a_8010_16807# distortionUnit_6.OUT a_7752_16807# VGND.t251 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X499 distortionUnit_5.tgate_1.IN distortionUnit_5.myOpamp_0.INn a_8134_23853# VGND.t91 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X500 a_20934_16677# a_20934_16677# VPWR.t166 VPWR.t165 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X501 a_8134_23853# a_7032_23398# VGND.t145 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X502 VPWR.t14 a_7876_23853# a_7876_23853# VPWR.t13 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X503 distortionUnit_3.tgate_1.IN ui_in[2].t19 distortionUnit_4.IN VGND.t32 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X504 VGND.t211 VGND.t210 VGND.t211 VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X505 bufferUnit_0.tgate_1.IN a_7736_36483# VPWR.t209 VPWR.t208 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X506 VGND.t209 VGND.t206 VGND.t208 VGND.t207 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0 ps=0 w=0.42 l=1
X507 VPWR.t136 ui_in[5].t19 distortionUnit_6.tgate_1.CTRLB distortionUnit_6.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X508 a_7876_23853# distortionUnit_5.IN.t16 a_8134_23853# VGND.t38 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X509 VPWR a_6912_30102# VGND sky130_fd_pr__res_xhigh_po_0p35 l=26.11
R0 ui_in[4].n2 ui_in[4].t9 212.081
R1 ui_in[4].n1 ui_in[4].t13 212.081
R2 ui_in[4].n6 ui_in[4].t15 212.081
R3 ui_in[4].n0 ui_in[4].t8 212.081
R4 ui_in[4].n11 ui_in[4].t10 212.081
R5 ui_in[4].n17 ui_in[4].t7 212.081
R6 ui_in[4].n12 ui_in[4].t5 212.081
R7 ui_in[4].n13 ui_in[4].t14 212.081
R8 ui_in[4] ui_in[4].n14 163.264
R9 ui_in[4].n16 ui_in[4].n15 152
R10 ui_in[4].n19 ui_in[4].n18 152
R11 ui_in[4].n10 ui_in[4].n9 152
R12 ui_in[4].n8 ui_in[4].n7 152
R13 ui_in[4].n5 ui_in[4].n4 152
R14 ui_in[4] ui_in[4].n3 152
R15 ui_in[4].n2 ui_in[4].t19 139.78
R16 ui_in[4].n1 ui_in[4].t2 139.78
R17 ui_in[4].n6 ui_in[4].t4 139.78
R18 ui_in[4].n0 ui_in[4].t18 139.78
R19 ui_in[4].n11 ui_in[4].t0 139.78
R20 ui_in[4].n17 ui_in[4].t17 139.78
R21 ui_in[4].n12 ui_in[4].t11 139.78
R22 ui_in[4].n13 ui_in[4].t3 139.78
R23 ui_in[4].n24 ui_in[4].t16 120.23
R24 ui_in[4].n24 ui_in[4].t6 120.228
R25 ui_in[4].n21 ui_in[4].t1 118.061
R26 ui_in[4].n21 ui_in[4].t12 118.058
R27 ui_in[4].n3 ui_in[4].n2 30.6732
R28 ui_in[4].n3 ui_in[4].n1 30.6732
R29 ui_in[4].n5 ui_in[4].n1 30.6732
R30 ui_in[4].n6 ui_in[4].n5 30.6732
R31 ui_in[4].n7 ui_in[4].n6 30.6732
R32 ui_in[4].n7 ui_in[4].n0 30.6732
R33 ui_in[4].n10 ui_in[4].n0 30.6732
R34 ui_in[4].n11 ui_in[4].n10 30.6732
R35 ui_in[4].n18 ui_in[4].n11 30.6732
R36 ui_in[4].n18 ui_in[4].n17 30.6732
R37 ui_in[4].n17 ui_in[4].n16 30.6732
R38 ui_in[4].n16 ui_in[4].n12 30.6732
R39 ui_in[4].n14 ui_in[4].n12 30.6732
R40 ui_in[4].n14 ui_in[4].n13 30.6732
R41 ui_in[4].n4 ui_in[4] 21.5045
R42 ui_in[4].n8 ui_in[4] 19.4565
R43 ui_in[4].n9 ui_in[4] 17.4085
R44 ui_in[4].n15 ui_in[4] 13.3125
R45 ui_in[4].n20 ui_in[4].n19 13.0565
R46 ui_in[4].n15 ui_in[4] 10.2405
R47 ui_in[4].n19 ui_in[4] 8.1925
R48 ui_in[4].n9 ui_in[4] 6.1445
R49 ui_in[4] ui_in[4].n8 4.0965
R50 ui_in[4].n23 ui_in[4].n20 3.2054
R51 ui_in[4].n20 ui_in[4] 2.3045
R52 ui_in[4].n4 ui_in[4] 2.0485
R53 ui_in[4].n22 ui_in[4].n21 0.528909
R54 ui_in[4].n25 ui_in[4].n24 0.506182
R55 ui_in[4].n26 ui_in[4].n25 0.42675
R56 ui_in[4].n26 ui_in[4].n23 0.342556
R57 ui_in[4].n23 ui_in[4].n22 0.3415
R58 ui_in[4].n25 ui_in[4] 0.170955
R59 ui_in[4].n22 ui_in[4] 0.148227
R60 ui_in[4] ui_in[4].n26 0.01225
R61 VGND.n551 VGND.n550 796000
R62 VGND.n537 VGND.n75 734302
R63 VGND.n538 VGND.n537 494301
R64 VGND.n1016 VGND.n543 488258
R65 VGND.n605 VGND.n543 405746
R66 VGND.n1045 VGND.n52 398767
R67 VGND.n1020 VGND.n1019 397063
R68 VGND.n1009 VGND.n551 324800
R69 VGND.n1009 VGND.n1008 284230
R70 VGND.n261 VGND.n150 137195
R71 VGND.n550 VGND.n549 122196
R72 VGND.n362 VGND.n335 98572.6
R73 VGND.n262 VGND 82857.8
R74 VGND.n725 VGND.n582 54678.4
R75 VGND.n153 VGND.n150 41031.3
R76 VGND.n153 VGND.n152 39882.8
R77 VGND.n230 VGND.n229 27500
R78 VGND.n481 VGND.n474 27500
R79 VGND.n710 VGND.n703 27500
R80 VGND.n793 VGND.n792 27500
R81 VGND.n994 VGND.n987 27500
R82 VGND.n931 VGND.n924 27500
R83 VGND.n304 VGND.n303 27500
R84 VGND.n426 VGND.n419 27500
R85 VGND.n827 VGND.n582 19915.8
R86 VGND.n828 VGND.n827 19476.5
R87 VGND.n262 VGND.n261 14154.2
R88 VGND.n230 VGND.t72 10325.8
R89 VGND.t51 VGND.n481 10325.8
R90 VGND.t193 VGND.n710 10325.8
R91 VGND.n793 VGND.t194 10325.8
R92 VGND.t152 VGND.n994 10325.8
R93 VGND.t195 VGND.n931 10325.8
R94 VGND.n304 VGND.t448 10325.8
R95 VGND.t382 VGND.n426 10325.8
R96 VGND.n242 VGND.n224 10285.8
R97 VGND.n483 VGND.n442 10285.8
R98 VGND.n712 VGND.n685 10285.8
R99 VGND.n805 VGND.n787 10285.8
R100 VGND.n996 VGND.n955 10285.8
R101 VGND.n933 VGND.n892 10285.8
R102 VGND.n316 VGND.n298 10285.8
R103 VGND.n428 VGND.n387 10285.8
R104 VGND.n231 VGND.n224 10253
R105 VGND.n480 VGND.n442 10253
R106 VGND.n709 VGND.n685 10253
R107 VGND.n794 VGND.n787 10253
R108 VGND.n993 VGND.n955 10253
R109 VGND.n930 VGND.n892 10253
R110 VGND.n305 VGND.n298 10253
R111 VGND.n425 VGND.n387 10253
R112 VGND.n242 VGND.n225 10250
R113 VGND.n483 VGND.n443 10250
R114 VGND.n712 VGND.n686 10250
R115 VGND.n805 VGND.n788 10250
R116 VGND.n996 VGND.n956 10250
R117 VGND.n933 VGND.n893 10250
R118 VGND.n316 VGND.n299 10250
R119 VGND.n428 VGND.n388 10250
R120 VGND.n231 VGND.n225 10187.3
R121 VGND.n480 VGND.n443 10187.3
R122 VGND.n709 VGND.n686 10187.3
R123 VGND.n794 VGND.n788 10187.3
R124 VGND.n993 VGND.n956 10187.3
R125 VGND.n930 VGND.n893 10187.3
R126 VGND.n305 VGND.n299 10187.3
R127 VGND.n425 VGND.n388 10187.3
R128 VGND.n942 VGND.n67 9815.24
R129 VGND.n1027 VGND.n67 9815.24
R130 VGND.n1027 VGND.n68 9815.24
R131 VGND.n160 VGND.n155 9815.24
R132 VGND.n257 VGND.n155 9815.24
R133 VGND.n257 VGND.n156 9815.24
R134 VGND.n87 VGND.n83 9815.24
R135 VGND.n529 VGND.n83 9815.24
R136 VGND.n529 VGND.n89 9815.24
R137 VGND.n592 VGND.n585 9815.24
R138 VGND.n824 VGND.n585 9815.24
R139 VGND.n824 VGND.n586 9815.24
R140 VGND.n49 VGND.n36 9815.24
R141 VGND.n1054 VGND.n36 9815.24
R142 VGND.n1054 VGND.n37 9815.24
R143 VGND.n134 VGND.n129 9815.24
R144 VGND.n331 VGND.n129 9815.24
R145 VGND.n331 VGND.n130 9815.24
R146 VGND.n368 VGND.n364 9815.24
R147 VGND.n373 VGND.n364 9815.24
R148 VGND.n373 VGND.n365 9815.24
R149 VGND.n1011 VGND.n548 8183.45
R150 VGND.n1016 VGND.n1015 8041.78
R151 VGND.n726 VGND.n725 6870.18
R152 VGND.n358 VGND.n337 6732.76
R153 VGND.n340 VGND.n339 6732.76
R154 VGND.n1040 VGND.n56 6732.76
R155 VGND.n61 VGND.n60 6732.76
R156 VGND.n753 VGND.n722 6732.76
R157 VGND.n600 VGND.n596 6732.76
R158 VGND.n609 VGND.n604 6732.76
R159 VGND.n558 VGND.n557 6732.76
R160 VGND.n1007 VGND.n552 6732.76
R161 VGND.n734 VGND.n728 6732.76
R162 VGND.n831 VGND.n569 6732.76
R163 VGND.n576 VGND.n571 6732.76
R164 VGND.n148 VGND.n142 6732.76
R165 VGND.n521 VGND.n92 6732.76
R166 VGND.n1061 VGND.n30 6732.76
R167 VGND.n539 VGND.n538 6359.87
R168 VGND.n526 VGND.n76 6338.76
R169 VGND.n535 VGND.n76 6338.76
R170 VGND.n526 VGND.n77 6338.76
R171 VGND.n535 VGND.n77 6338.76
R172 VGND.n1023 VGND.n72 6338.76
R173 VGND.n73 VGND.n72 6338.76
R174 VGND.n1023 VGND.n1022 6338.76
R175 VGND.n1022 VGND.n73 6338.76
R176 VGND.n251 VGND.n166 6338.76
R177 VGND.n251 VGND.n167 6338.76
R178 VGND.n252 VGND.n166 6338.76
R179 VGND.n252 VGND.n167 6338.76
R180 VGND.n815 VGND.n813 6338.76
R181 VGND.n817 VGND.n813 6338.76
R182 VGND.n816 VGND.n815 6338.76
R183 VGND.n817 VGND.n816 6338.76
R184 VGND.n46 VGND.n44 6338.76
R185 VGND.n1047 VGND.n44 6338.76
R186 VGND.n47 VGND.n46 6338.76
R187 VGND.n1047 VGND.n47 6338.76
R188 VGND.n325 VGND.n140 6338.76
R189 VGND.n325 VGND.n141 6338.76
R190 VGND.n326 VGND.n140 6338.76
R191 VGND.n326 VGND.n141 6338.76
R192 VGND.n376 VGND.n127 6338.76
R193 VGND.n376 VGND.n124 6338.76
R194 VGND.n377 VGND.n127 6338.76
R195 VGND.n377 VGND.n124 6338.76
R196 VGND.n1017 VGND.n539 5925.42
R197 VGND.n1014 VGND.n545 5515.01
R198 VGND.n1045 VGND.n1044 5420.28
R199 VGND.n605 VGND.n544 4759.63
R200 VGND.n538 VGND.n74 4034.2
R201 VGND.n1020 VGND.n539 3806.52
R202 VGND.n1044 VGND.n53 3806.09
R203 VGND.n741 VGND.n545 3676.5
R204 VGND.n267 VGND.n266 3671.5
R205 VGND.n1043 VGND.n1042 3434.11
R206 VGND.n338 VGND.n337 3366.38
R207 VGND.n350 VGND.n339 3366.38
R208 VGND.n1040 VGND.n57 3366.38
R209 VGND.n1033 VGND.n60 3366.38
R210 VGND.n753 VGND.n723 3366.38
R211 VGND.n600 VGND.n599 3366.38
R212 VGND.n609 VGND.n608 3366.38
R213 VGND.n562 VGND.n557 3366.38
R214 VGND.n1007 VGND.n555 3366.38
R215 VGND.n734 VGND.n731 3366.38
R216 VGND.n831 VGND.n570 3366.38
R217 VGND.n576 VGND.n573 3366.38
R218 VGND.n145 VGND.n142 3366.38
R219 VGND.n521 VGND.n93 3366.38
R220 VGND.n1061 VGND.n31 3366.38
R221 VGND.n65 VGND.n54 3016.93
R222 VGND.n1010 VGND.n550 3001.37
R223 VGND.n724 VGND 2969.99
R224 VGND.n1015 VGND.n1014 2508.09
R225 VGND.n345 VGND.n344 2399.08
R226 VGND.n580 VGND.n578 2198.58
R227 VGND.n344 VGND.n32 2191.03
R228 VGND.n266 VGND.n91 2083.37
R229 VGND.n581 VGND.n580 2036.22
R230 VGND.n737 VGND.n736 1920.23
R231 VGND.n524 VGND.n90 1850.51
R232 VGND.n362 VGND.n361 1822.86
R233 VGND.n738 VGND.n737 1776.8
R234 VGND.n742 VGND.n739 1683.19
R235 VGND.n747 VGND.n739 1683.19
R236 VGND.n1015 VGND.n544 1504.19
R237 VGND.n1017 VGND.n1016 1483.43
R238 VGND.n347 VGND.n346 1478.96
R239 VGND.n265 VGND.n53 1460.08
R240 VGND.n1013 VGND.n1012 1386.21
R241 VGND.n347 VGND.n345 1330.05
R242 VGND.n229 VGND.t242 1302.55
R243 VGND.n474 VGND.t332 1302.55
R244 VGND.n703 VGND.t222 1302.55
R245 VGND.n792 VGND.t261 1302.55
R246 VGND.n987 VGND.t288 1302.55
R247 VGND.n924 VGND.t233 1302.55
R248 VGND.n303 VGND.t245 1302.55
R249 VGND.n419 VGND.t282 1302.55
R250 VGND.n523 VGND.n91 1281.68
R251 VGND.n578 VGND.n32 1243.6
R252 VGND.n1057 VGND.n1056 1234.1
R253 VGND.n749 VGND.n545 1234.1
R254 VGND.n1030 VGND.n1029 1234.1
R255 VGND.n1018 VGND.n541 1234.1
R256 VGND.t386 VGND.n584 1231.2
R257 VGND.t386 VGND.n548 1231.2
R258 VGND.n741 VGND.n738 1229.9
R259 VGND.n736 VGND.n581 1221.82
R260 VGND.n1041 VGND.t78 1198.65
R261 VGND.n63 VGND.t79 1198.65
R262 VGND.t119 VGND.n546 1198.65
R263 VGND.t118 VGND.n597 1198.65
R264 VGND.t456 VGND.n559 1198.65
R265 VGND.t455 VGND.n560 1198.65
R266 VGND.n735 VGND.t421 1198.65
R267 VGND.t420 VGND.n729 1198.65
R268 VGND.t171 VGND.n743 1198.65
R269 VGND.n748 VGND.t170 1198.65
R270 VGND.n577 VGND.t86 1198.65
R271 VGND.t87 VGND.n33 1198.65
R272 VGND.t392 VGND.n143 1198.65
R273 VGND.n149 VGND.t393 1198.65
R274 VGND.n342 VGND.t458 1198.65
R275 VGND.n359 VGND.t457 1198.65
R276 VGND.n259 VGND.n153 1160.48
R277 VGND.n1010 VGND.n1009 1124.01
R278 VGND.n1009 VGND.n54 1124.01
R279 VGND.n827 VGND.n826 1083.35
R280 VGND.n333 VGND.n34 1063.33
R281 VGND.n589 VGND.n583 1063.33
R282 VGND.n260 VGND.n64 1063.33
R283 VGND.t59 VGND.n66 1055.41
R284 VGND.t59 VGND.n1021 1055.41
R285 VGND.t15 VGND.n55 1053.4
R286 VGND.t6 VGND.n1031 1053.4
R287 VGND.n752 VGND.t426 1053.4
R288 VGND.t18 VGND.n750 1053.4
R289 VGND.t174 VGND.n547 1053.4
R290 VGND.t122 VGND.n606 1053.4
R291 VGND.n1008 VGND.t31 1053.4
R292 VGND.t32 VGND.n553 1053.4
R293 VGND.n830 VGND.t33 1053.4
R294 VGND.t163 VGND.n828 1053.4
R295 VGND.n522 VGND.t65 1053.4
R296 VGND.n152 VGND.t427 1053.4
R297 VGND.t139 VGND.n348 1053.4
R298 VGND.t109 VGND.n336 1053.4
R299 VGND.n1060 VGND.t52 1053.4
R300 VGND.t140 VGND.n1058 1053.4
R301 VGND.t62 VGND.n35 1040.9
R302 VGND.n1046 VGND.t62 1040.9
R303 VGND.t469 VGND.n128 962.694
R304 VGND.t469 VGND.n267 962.694
R305 VGND.t88 VGND.n154 962.694
R306 VGND.t88 VGND.n74 962.694
R307 VGND.n1018 VGND.n1017 957.76
R308 VGND.n745 VGND.n739 841.596
R309 VGND.t242 VGND.t91 803.966
R310 VGND.t91 VGND.t36 803.966
R311 VGND.t36 VGND.t146 803.966
R312 VGND.t146 VGND.t95 803.966
R313 VGND.t95 VGND.t94 803.966
R314 VGND.t37 VGND.t38 803.966
R315 VGND.t93 VGND.t92 803.966
R316 VGND.t236 VGND.t93 803.966
R317 VGND.t301 VGND.t236 803.966
R318 VGND.t332 VGND.t358 803.966
R319 VGND.t358 VGND.t251 803.966
R320 VGND.t251 VGND.t101 803.966
R321 VGND.t101 VGND.t103 803.966
R322 VGND.t103 VGND.t105 803.966
R323 VGND.t107 VGND.t99 803.966
R324 VGND.t97 VGND.t298 803.966
R325 VGND.t298 VGND.t309 803.966
R326 VGND.t309 VGND.t323 803.966
R327 VGND.t222 VGND.t213 803.966
R328 VGND.t213 VGND.t293 803.966
R329 VGND.t293 VGND.t96 803.966
R330 VGND.t96 VGND.t418 803.966
R331 VGND.t418 VGND.t411 803.966
R332 VGND.t409 VGND.t413 803.966
R333 VGND.t415 VGND.t363 803.966
R334 VGND.t363 VGND.t219 803.966
R335 VGND.t219 VGND.t207 803.966
R336 VGND.t261 VGND.t279 803.966
R337 VGND.t279 VGND.t326 803.966
R338 VGND.t326 VGND.t446 803.966
R339 VGND.t446 VGND.t408 803.966
R340 VGND.t408 VGND.t406 803.966
R341 VGND.t440 VGND.t443 803.966
R342 VGND.t377 VGND.t407 803.966
R343 VGND.t264 VGND.t377 803.966
R344 VGND.t216 VGND.t264 803.966
R345 VGND.t288 VGND.t276 803.966
R346 VGND.t276 VGND.t74 803.966
R347 VGND.t74 VGND.t75 803.966
R348 VGND.t75 VGND.t381 803.966
R349 VGND.t381 VGND.t380 803.966
R350 VGND.t77 VGND.t73 803.966
R351 VGND.t379 VGND.t239 803.966
R352 VGND.t239 VGND.t76 803.966
R353 VGND.t76 VGND.t267 803.966
R354 VGND.t233 VGND.t346 803.966
R355 VGND.t346 VGND.t42 803.966
R356 VGND.t42 VGND.t43 803.966
R357 VGND.t43 VGND.t159 803.966
R358 VGND.t159 VGND.t157 803.966
R359 VGND.t40 VGND.t41 803.966
R360 VGND.t154 VGND.t227 803.966
R361 VGND.t227 VGND.t44 803.966
R362 VGND.t44 VGND.t248 803.966
R363 VGND.t245 VGND.t285 803.966
R364 VGND.t285 VGND.t273 803.966
R365 VGND.t273 VGND.t190 803.966
R366 VGND.t190 VGND.t182 803.966
R367 VGND.t182 VGND.t180 803.966
R368 VGND.t186 VGND.t184 803.966
R369 VGND.t329 VGND.t188 803.966
R370 VGND.t370 VGND.t329 803.966
R371 VGND.t257 VGND.t370 803.966
R372 VGND.t282 VGND.t198 803.966
R373 VGND.t198 VGND.t204 803.966
R374 VGND.t204 VGND.t205 803.966
R375 VGND.t205 VGND.t196 803.966
R376 VGND.t196 VGND.t197 803.966
R377 VGND.t202 VGND.t203 803.966
R378 VGND.t199 VGND.t200 803.966
R379 VGND.t200 VGND.t201 803.966
R380 VGND.t201 VGND.t230 803.966
R381 VGND.n725 VGND.n583 795.182
R382 VGND.n537 VGND.n536 783.655
R383 VGND.n525 VGND.n524 774.306
R384 VGND.n524 VGND.n523 698.878
R385 VGND.n235 VGND.n226 666.376
R386 VGND.n485 VGND.n440 666.376
R387 VGND.n714 VGND.n683 666.376
R388 VGND.n798 VGND.n789 666.376
R389 VGND.n998 VGND.n953 666.376
R390 VGND.n935 VGND.n890 666.376
R391 VGND.n309 VGND.n300 666.376
R392 VGND.n430 VGND.n385 666.376
R393 VGND.n241 VGND.n240 665.019
R394 VGND.n484 VGND.n441 665.019
R395 VGND.n713 VGND.n684 665.019
R396 VGND.n804 VGND.n803 665.019
R397 VGND.n997 VGND.n954 665.019
R398 VGND.n934 VGND.n891 665.019
R399 VGND.n315 VGND.n314 665.019
R400 VGND.n429 VGND.n386 665.019
R401 VGND.n234 VGND.n233 664.242
R402 VGND.n477 VGND.n475 664.242
R403 VGND.n706 VGND.n704 664.242
R404 VGND.n797 VGND.n796 664.242
R405 VGND.n990 VGND.n988 664.242
R406 VGND.n927 VGND.n925 664.242
R407 VGND.n308 VGND.n307 664.242
R408 VGND.n422 VGND.n420 664.242
R409 VGND.n232 VGND.n227 661.915
R410 VGND.n479 VGND.n478 661.915
R411 VGND.n708 VGND.n707 661.915
R412 VGND.n795 VGND.n790 661.915
R413 VGND.n992 VGND.n991 661.915
R414 VGND.n929 VGND.n928 661.915
R415 VGND.n306 VGND.n301 661.915
R416 VGND.n424 VGND.n423 661.915
R417 VGND.n264 VGND.n263 660.718
R418 VGND.t72 VGND.t301 660.674
R419 VGND.t323 VGND.t51 660.674
R420 VGND.t207 VGND.t193 660.674
R421 VGND.t194 VGND.t216 660.674
R422 VGND.t267 VGND.t152 660.674
R423 VGND.t248 VGND.t195 660.674
R424 VGND.t448 VGND.t257 660.674
R425 VGND.t230 VGND.t382 660.674
R426 VGND.n263 VGND.n53 660.265
R427 VGND.n1026 VGND.n69 646.878
R428 VGND.n256 VGND.n157 637.741
R429 VGND.n161 VGND.n157 637.741
R430 VGND.n162 VGND.n161 637.741
R431 VGND.n86 VGND.n82 637.741
R432 VGND.n86 VGND.n84 637.741
R433 VGND.n530 VGND.n82 637.741
R434 VGND.n594 VGND.n593 637.741
R435 VGND.n593 VGND.n587 637.741
R436 VGND.n823 VGND.n587 637.741
R437 VGND.n944 VGND.n943 637.741
R438 VGND.n943 VGND.n69 637.741
R439 VGND.n48 VGND.n40 637.741
R440 VGND.n48 VGND.n38 637.741
R441 VGND.n1053 VGND.n38 637.741
R442 VGND.n330 VGND.n131 637.741
R443 VGND.n135 VGND.n131 637.741
R444 VGND.n136 VGND.n135 637.741
R445 VGND.n370 VGND.n369 637.741
R446 VGND.n369 VGND.n366 637.741
R447 VGND.n372 VGND.n370 637.741
R448 VGND.n62 VGND.t78 636.323
R449 VGND.t79 VGND.n62 636.323
R450 VGND.n598 VGND.t119 636.323
R451 VGND.n598 VGND.t118 636.323
R452 VGND.n561 VGND.t456 636.323
R453 VGND.n561 VGND.t455 636.323
R454 VGND.n730 VGND.t421 636.323
R455 VGND.n730 VGND.t420 636.323
R456 VGND.n744 VGND.t171 636.323
R457 VGND.n744 VGND.t170 636.323
R458 VGND.n572 VGND.t86 636.323
R459 VGND.n572 VGND.t87 636.323
R460 VGND.n144 VGND.t392 636.323
R461 VGND.n144 VGND.t393 636.323
R462 VGND.t458 VGND.n341 636.323
R463 VGND.n341 VGND.t457 636.323
R464 VGND.t38 VGND.n243 629.462
R465 VGND.n482 VGND.t99 629.462
R466 VGND.n711 VGND.t413 629.462
R467 VGND.t443 VGND.n806 629.462
R468 VGND.n995 VGND.t73 629.462
R469 VGND.n932 VGND.t41 629.462
R470 VGND.t184 VGND.n317 629.462
R471 VGND.n427 VGND.t203 629.462
R472 VGND.n261 VGND.n260 621.763
R473 VGND VGND.n542 620.966
R474 VGND.n525 VGND 581.288
R475 VGND.n346 VGND 581.236
R476 VGND.n343 VGND 562.322
R477 VGND.n579 VGND 560.347
R478 VGND.n65 VGND 559.942
R479 VGND.n1032 VGND.t15 559.212
R480 VGND.n1032 VGND.t6 559.212
R481 VGND.t426 VGND.n751 559.212
R482 VGND.n751 VGND.t18 559.212
R483 VGND.n607 VGND.t174 559.212
R484 VGND.n607 VGND.t122 559.212
R485 VGND.n554 VGND.t31 559.212
R486 VGND.n554 VGND.t32 559.212
R487 VGND.t33 VGND.n829 559.212
R488 VGND.n829 VGND.t163 559.212
R489 VGND.n151 VGND.t65 559.212
R490 VGND.t427 VGND.n151 559.212
R491 VGND.n349 VGND.t139 559.212
R492 VGND.n349 VGND.t109 559.212
R493 VGND.t52 VGND.n1059 559.212
R494 VGND.n1059 VGND.t140 559.212
R495 VGND.n727 VGND 554.649
R496 VGND.n549 VGND 552.415
R497 VGND.n1014 VGND.n1013 545.561
R498 VGND.n1056 VGND 524.37
R499 VGND.n1029 VGND.n1028 508.959
R500 VGND.n1029 VGND 504.416
R501 VGND.n1056 VGND.n1055 475.07
R502 VGND.n1012 VGND.n1011 461.769
R503 VGND.n1046 VGND.n1045 442.577
R504 VGND.n1021 VGND.n1020 435.115
R505 VGND.n1025 VGND.n70 432.467
R506 VGND.n825 VGND.n584 429.399
R507 VGND.n244 VGND.t94 414.449
R508 VGND.t105 VGND.n473 414.449
R509 VGND.t411 VGND.n702 414.449
R510 VGND.n807 VGND.t406 414.449
R511 VGND.t380 VGND.n986 414.449
R512 VGND.t157 VGND.n923 414.449
R513 VGND.n318 VGND.t180 414.449
R514 VGND.t197 VGND.n418 414.449
R515 VGND.n253 VGND.n165 411.495
R516 VGND.n534 VGND.n533 411.495
R517 VGND.n818 VGND.n812 411.495
R518 VGND.n1048 VGND.n43 411.495
R519 VGND.n327 VGND.n139 411.495
R520 VGND.n379 VGND.n378 411.495
R521 VGND.n947 VGND.n70 411.156
R522 VGND.n254 VGND.n253 398.683
R523 VGND.n533 VGND.n532 398.683
R524 VGND.n812 VGND.n588 398.683
R525 VGND.n43 VGND.n39 398.683
R526 VGND.n328 VGND.n327 398.683
R527 VGND.n378 VGND.n125 398.683
R528 VGND.n244 VGND.t37 389.519
R529 VGND.n473 VGND.t107 389.519
R530 VGND.n702 VGND.t409 389.519
R531 VGND.n807 VGND.t440 389.519
R532 VGND.n986 VGND.t77 389.519
R533 VGND.n923 VGND.t40 389.519
R534 VGND.n318 VGND.t186 389.519
R535 VGND.n418 VGND.t202 389.519
R536 VGND.n1028 VGND.n66 368.087
R537 VGND.n1055 VGND.n35 363.026
R538 VGND.n250 VGND.n164 347.647
R539 VGND.n324 VGND.n138 347.647
R540 VGND.n126 VGND.n123 347.647
R541 VGND.n80 VGND.n79 347.646
R542 VGND.n814 VGND.n811 347.646
R543 VGND.n45 VGND.n42 347.646
R544 VGND.n549 VGND.t68 343.673
R545 VGND.n332 VGND.n128 335.752
R546 VGND.n258 VGND.n154 335.752
R547 VGND.n727 VGND.t472 319.978
R548 VGND.n133 VGND.n130 315.68
R549 VGND.n50 VGND.n37 315.68
R550 VGND.n591 VGND.n586 315.68
R551 VGND.n89 VGND.n88 315.68
R552 VGND.n159 VGND.n156 315.68
R553 VGND.n941 VGND.n68 315.68
R554 VGND.n946 VGND.n71 300.587
R555 VGND.n531 VGND.n81 287.356
R556 VGND.n822 VGND.n821 287.356
R557 VGND.n1052 VGND.n1051 287.356
R558 VGND.n371 VGND.n122 287.356
R559 VGND.n255 VGND.n163 287.356
R560 VGND.n329 VGND.n137 287.356
R561 VGND.n182 VGND.t12 287.151
R562 VGND.n110 VGND.t111 287.151
R563 VGND.n655 VGND.t425 287.151
R564 VGND.n849 VGND.t454 287.151
R565 VGND.n505 VGND.t67 287.151
R566 VGND.n16 VGND.t56 287.151
R567 VGND.n367 VGND.n365 285.233
R568 VGND.n171 VGND.t1 284.024
R569 VGND.n99 VGND.t128 284.024
R570 VGND.n644 VGND.t473 284.024
R571 VGND.n838 VGND.t169 284.024
R572 VGND.n494 VGND.t431 284.024
R573 VGND.n5 VGND.t403 284.024
R574 VGND.n629 VGND.t178 282.885
R575 VGND.n876 VGND.t25 282.885
R576 VGND.n617 VGND.t69 280.457
R577 VGND.n864 VGND.t83 280.457
R578 VGND.n266 VGND.n265 278.738
R579 VGND.t438 VGND.n132 277.17
R580 VGND.n51 VGND.t153 277.17
R581 VGND.t39 VGND.n590 277.17
R582 VGND.t23 VGND.n85 277.17
R583 VGND.t192 VGND.n158 277.17
R584 VGND.t179 VGND.n540 277.17
R585 VGND.n826 VGND.n825 274.337
R586 VGND.t389 VGND.n375 265.567
R587 VGND.t389 VGND.n90 265.567
R588 VGND.t82 VGND.n65 265.002
R589 VGND.n527 VGND.t383 263.87
R590 VGND.n536 VGND.t383 263.87
R591 VGND.n1042 VGND.n1041 261.435
R592 VGND.n1030 VGND.n63 261.435
R593 VGND.n1013 VGND.n546 261.435
R594 VGND.n597 VGND.n544 261.435
R595 VGND.n559 VGND.n551 261.435
R596 VGND.n560 VGND.n541 261.435
R597 VGND.n736 VGND.n735 261.435
R598 VGND.n729 VGND.n582 261.435
R599 VGND.n743 VGND.n741 261.435
R600 VGND.n749 VGND.n748 261.435
R601 VGND.n578 VGND.n577 261.435
R602 VGND.n1057 VGND.n33 261.435
R603 VGND.n143 VGND.n91 261.435
R604 VGND.n150 VGND.n149 261.435
R605 VGND.n345 VGND.n342 261.435
R606 VGND.n360 VGND.n359 261.435
R607 VGND.n579 VGND.t168 260.86
R608 VGND.n263 VGND 257.546
R609 VGND.n945 VGND.n71 255.356
R610 VGND.n747 VGND.n746 254.685
R611 VGND.n528 VGND 253.361
R612 VGND.n343 VGND.t402 240.785
R613 VGND.n216 VGND.t303 236.113
R614 VGND.n464 VGND.t354 236.113
R615 VGND.n693 VGND.t209 236.113
R616 VGND.n779 VGND.t255 236.113
R617 VGND.n977 VGND.t269 236.113
R618 VGND.n914 VGND.t336 236.113
R619 VGND.n290 VGND.t259 236.113
R620 VGND.n409 VGND.t317 236.113
R621 VGND.t243 VGND.n200 235.764
R622 VGND.t366 VGND.n447 235.764
R623 VGND.t223 VGND.n670 235.764
R624 VGND.t307 VGND.n763 235.764
R625 VGND.t289 VGND.n960 235.764
R626 VGND.t319 VGND.n897 235.764
R627 VGND.t246 VGND.n274 235.764
R628 VGND.t351 VGND.n392 235.764
R629 VGND.n333 VGND.n332 233.161
R630 VGND.n358 VGND.n357 232.597
R631 VGND.n351 VGND.n340 232.597
R632 VGND.n58 VGND.n56 232.597
R633 VGND.n1034 VGND.n61 232.597
R634 VGND.n722 VGND.n721 232.597
R635 VGND.n596 VGND.n595 232.597
R636 VGND.n604 VGND.n603 232.597
R637 VGND.n563 VGND.n558 232.597
R638 VGND.n556 VGND.n552 232.597
R639 VGND.n732 VGND.n728 232.597
R640 VGND.n569 VGND.n568 232.597
R641 VGND.n574 VGND.n571 232.597
R642 VGND.n148 VGND.n147 232.597
R643 VGND.n94 VGND.n92 232.597
R644 VGND.n30 VGND.n29 232.597
R645 VGND.n1042 VGND.n55 229.755
R646 VGND.n1031 VGND.n1030 229.755
R647 VGND.n752 VGND.n738 229.755
R648 VGND.n750 VGND.n749 229.755
R649 VGND.n1012 VGND.n547 229.755
R650 VGND.n606 VGND.n605 229.755
R651 VGND.n553 VGND.n541 229.755
R652 VGND.n830 VGND.n581 229.755
R653 VGND.n523 VGND.n522 229.755
R654 VGND.n348 VGND.n347 229.755
R655 VGND.n360 VGND.n336 229.755
R656 VGND.n1060 VGND.n32 229.755
R657 VGND.n1058 VGND.n1057 229.755
R658 VGND VGND.n335 220.334
R659 VGND.n176 VGND.n170 207.213
R660 VGND.n189 VGND.n177 207.213
R661 VGND.n179 VGND.n178 207.213
R662 VGND.n104 VGND.n98 207.213
R663 VGND.n117 VGND.n105 207.213
R664 VGND.n107 VGND.n106 207.213
R665 VGND.n623 VGND.n616 207.213
R666 VGND.n636 VGND.n624 207.213
R667 VGND.n626 VGND.n625 207.213
R668 VGND.n649 VGND.n643 207.213
R669 VGND.n662 VGND.n650 207.213
R670 VGND.n652 VGND.n651 207.213
R671 VGND.n870 VGND.n863 207.213
R672 VGND.n883 VGND.n871 207.213
R673 VGND.n873 VGND.n872 207.213
R674 VGND.n843 VGND.n837 207.213
R675 VGND.n856 VGND.n844 207.213
R676 VGND.n846 VGND.n845 207.213
R677 VGND.n499 VGND.n493 207.213
R678 VGND.n512 VGND.n500 207.213
R679 VGND.n502 VGND.n501 207.213
R680 VGND.n10 VGND.n4 207.213
R681 VGND.n23 VGND.n11 207.213
R682 VGND.n13 VGND.n12 207.213
R683 VGND.n167 VGND.n165 199.829
R684 VGND.n535 VGND.n534 199.829
R685 VGND.n818 VGND.n817 199.829
R686 VGND.n947 VGND.n73 199.829
R687 VGND.n1048 VGND.n1047 199.829
R688 VGND.n141 VGND.n139 199.829
R689 VGND.n379 VGND.n124 199.829
R690 VGND.n124 VGND.n90 195
R691 VGND.n127 VGND.n126 195
R692 VGND.n375 VGND.n127 195
R693 VGND.n373 VGND.n372 195
R694 VGND.n374 VGND.n373 195
R695 VGND.n369 VGND.n368 195
R696 VGND.n267 VGND.n141 195
R697 VGND.n140 VGND.n138 195
R698 VGND.n140 VGND.n128 195
R699 VGND.n331 VGND.n330 195
R700 VGND.n332 VGND.n331 195
R701 VGND.n135 VGND.n134 195
R702 VGND.n1047 VGND.n1046 195
R703 VGND.n46 VGND.n45 195
R704 VGND.n46 VGND.n35 195
R705 VGND.n1054 VGND.n1053 195
R706 VGND.n1055 VGND.n1054 195
R707 VGND.n49 VGND.n48 195
R708 VGND.n817 VGND.n548 195
R709 VGND.n815 VGND.n814 195
R710 VGND.n815 VGND.n584 195
R711 VGND.n824 VGND.n823 195
R712 VGND.n825 VGND.n824 195
R713 VGND.n593 VGND.n592 195
R714 VGND.n87 VGND.n86 195
R715 VGND.n167 VGND.n74 195
R716 VGND.n166 VGND.n164 195
R717 VGND.n166 VGND.n154 195
R718 VGND.n257 VGND.n256 195
R719 VGND.n258 VGND.n257 195
R720 VGND.n161 VGND.n160 195
R721 VGND.n1021 VGND.n73 195
R722 VGND.n1024 VGND.n1023 195
R723 VGND.n1023 VGND.n66 195
R724 VGND.n1027 VGND.n1026 195
R725 VGND.n1028 VGND.n1027 195
R726 VGND.n943 VGND.n942 195
R727 VGND.n536 VGND.n535 195
R728 VGND.n526 VGND.n80 195
R729 VGND.n527 VGND.n526 195
R730 VGND.n530 VGND.n529 195
R731 VGND.n529 VGND.n528 195
R732 VGND.n221 VGND.n220 194.805
R733 VGND.n469 VGND.n468 194.805
R734 VGND.n698 VGND.n697 194.805
R735 VGND.n784 VGND.n783 194.805
R736 VGND.n982 VGND.n981 194.805
R737 VGND.n919 VGND.n918 194.805
R738 VGND.n295 VGND.n294 194.805
R739 VGND.n414 VGND.n413 194.805
R740 VGND.n207 VGND.n206 194.542
R741 VGND.n454 VGND.n453 194.542
R742 VGND.n677 VGND.n676 194.542
R743 VGND.n770 VGND.n769 194.542
R744 VGND.n967 VGND.n966 194.542
R745 VGND.n904 VGND.n903 194.542
R746 VGND.n281 VGND.n280 194.542
R747 VGND.n399 VGND.n398 194.542
R748 VGND.n223 VGND.n222 194.463
R749 VGND.n209 VGND.n208 194.463
R750 VGND.n471 VGND.n470 194.463
R751 VGND.n456 VGND.n455 194.463
R752 VGND.n700 VGND.n699 194.463
R753 VGND.n679 VGND.n678 194.463
R754 VGND.n786 VGND.n785 194.463
R755 VGND.n772 VGND.n771 194.463
R756 VGND.n984 VGND.n983 194.463
R757 VGND.n969 VGND.n968 194.463
R758 VGND.n921 VGND.n920 194.463
R759 VGND.n906 VGND.n905 194.463
R760 VGND.n297 VGND.n296 194.463
R761 VGND.n283 VGND.n282 194.463
R762 VGND.n416 VGND.n415 194.463
R763 VGND.n401 VGND.n400 194.463
R764 VGND.n217 VGND.n216 194.3
R765 VGND.n219 VGND.n218 194.3
R766 VGND.n205 VGND.n204 194.3
R767 VGND.n202 VGND.n201 194.3
R768 VGND.n465 VGND.n464 194.3
R769 VGND.n467 VGND.n466 194.3
R770 VGND.n452 VGND.n451 194.3
R771 VGND.n449 VGND.n448 194.3
R772 VGND.n694 VGND.n693 194.3
R773 VGND.n696 VGND.n695 194.3
R774 VGND.n675 VGND.n674 194.3
R775 VGND.n672 VGND.n671 194.3
R776 VGND.n780 VGND.n779 194.3
R777 VGND.n782 VGND.n781 194.3
R778 VGND.n768 VGND.n767 194.3
R779 VGND.n765 VGND.n764 194.3
R780 VGND.n978 VGND.n977 194.3
R781 VGND.n980 VGND.n979 194.3
R782 VGND.n965 VGND.n964 194.3
R783 VGND.n962 VGND.n961 194.3
R784 VGND.n915 VGND.n914 194.3
R785 VGND.n917 VGND.n916 194.3
R786 VGND.n902 VGND.n901 194.3
R787 VGND.n899 VGND.n898 194.3
R788 VGND.n291 VGND.n290 194.3
R789 VGND.n293 VGND.n292 194.3
R790 VGND.n279 VGND.n278 194.3
R791 VGND.n276 VGND.n275 194.3
R792 VGND.n410 VGND.n409 194.3
R793 VGND.n412 VGND.n411 194.3
R794 VGND.n397 VGND.n396 194.3
R795 VGND.n394 VGND.n393 194.3
R796 VGND.n264 VGND.t0 190.006
R797 VGND.n229 VGND.n224 189.166
R798 VGND.n474 VGND.n442 189.166
R799 VGND.n703 VGND.n685 189.166
R800 VGND.n792 VGND.n787 189.166
R801 VGND.n987 VGND.n955 189.166
R802 VGND.n924 VGND.n892 189.166
R803 VGND.n303 VGND.n298 189.166
R804 VGND.n419 VGND.n387 189.166
R805 VGND.n368 VGND.n367 185.647
R806 VGND.n942 VGND.n941 185.053
R807 VGND.n160 VGND.n159 185.053
R808 VGND.n88 VGND.n87 185.053
R809 VGND.n592 VGND.n591 185.053
R810 VGND.n50 VGND.n49 185.053
R811 VGND.n134 VGND.n133 185.053
R812 VGND.n363 VGND.n362 182.97
R813 VGND.n334 VGND.n333 181.347
R814 VGND.n1056 VGND.n34 180.559
R815 VGND.n589 VGND.n545 180.559
R816 VGND.n1029 VGND.n64 180.559
R817 VGND.n1019 VGND.n1018 180.559
R818 VGND.n243 VGND.t92 174.505
R819 VGND.n482 VGND.t97 174.505
R820 VGND.n711 VGND.t415 174.505
R821 VGND.n806 VGND.t407 174.505
R822 VGND.n995 VGND.t379 174.505
R823 VGND.n932 VGND.t154 174.505
R824 VGND.n317 VGND.t188 174.505
R825 VGND.n427 VGND.t199 174.505
R826 VGND.n259 VGND.n258 168.912
R827 VGND.n1017 VGND.n542 165.303
R828 VGND.n580 VGND.n579 163.56
R829 VGND.n344 VGND.n343 151.095
R830 VGND.n356 VGND.n337 147.038
R831 VGND.n1040 VGND.n1039 147.038
R832 VGND.n1035 VGND.n60 147.038
R833 VGND.n754 VGND.n753 147.038
R834 VGND.n601 VGND.n600 147.038
R835 VGND.n610 VGND.n609 147.038
R836 VGND.n564 VGND.n557 147.038
R837 VGND.n1007 VGND.n1006 147.038
R838 VGND.n734 VGND.n733 147.038
R839 VGND.n832 VGND.n831 147.038
R840 VGND.n742 VGND.n740 147.038
R841 VGND.n576 VGND.n575 147.038
R842 VGND.n146 VGND.n142 147.038
R843 VGND.n521 VGND.n520 147.038
R844 VGND.n352 VGND.n339 147.038
R845 VGND.n1062 VGND.n1061 147.038
R846 VGND.n1031 VGND.n61 146.25
R847 VGND.n60 VGND.n55 146.25
R848 VGND.n63 VGND.n56 146.25
R849 VGND.n1041 VGND.n1040 146.25
R850 VGND.n750 VGND.n722 146.25
R851 VGND.n753 VGND.n752 146.25
R852 VGND.n597 VGND.n596 146.25
R853 VGND.n600 VGND.n546 146.25
R854 VGND.n606 VGND.n604 146.25
R855 VGND.n609 VGND.n547 146.25
R856 VGND.n560 VGND.n558 146.25
R857 VGND.n559 VGND.n557 146.25
R858 VGND.n553 VGND.n552 146.25
R859 VGND.n1008 VGND.n1007 146.25
R860 VGND.n729 VGND.n728 146.25
R861 VGND.n735 VGND.n734 146.25
R862 VGND.n828 VGND.n569 146.25
R863 VGND.n831 VGND.n830 146.25
R864 VGND.n743 VGND.n742 146.25
R865 VGND.n748 VGND.n747 146.25
R866 VGND.n571 VGND.n33 146.25
R867 VGND.n577 VGND.n576 146.25
R868 VGND.n149 VGND.n148 146.25
R869 VGND.n143 VGND.n142 146.25
R870 VGND.n152 VGND.n92 146.25
R871 VGND.n522 VGND.n521 146.25
R872 VGND.n340 VGND.n336 146.25
R873 VGND.n348 VGND.n339 146.25
R874 VGND.n359 VGND.n358 146.25
R875 VGND.n342 VGND.n337 146.25
R876 VGND.n1058 VGND.n30 146.25
R877 VGND.n1061 VGND.n1060 146.25
R878 VGND.t68 VGND.t175 144.262
R879 VGND.t175 VGND.t120 144.262
R880 VGND.t120 VGND.t125 144.262
R881 VGND.t125 VGND.t70 144.262
R882 VGND.t70 VGND.t123 144.262
R883 VGND.t123 VGND.t172 144.262
R884 VGND.t472 VGND.t461 134.107
R885 VGND.t461 VGND.t21 134.107
R886 VGND.t21 VGND.t422 134.107
R887 VGND.t422 VGND.t459 134.107
R888 VGND.t459 VGND.t19 134.107
R889 VGND.t19 VGND.t474 134.107
R890 VGND.t474 VGND.n726 124.528
R891 VGND.n1043 VGND.n54 122.853
R892 VGND.n335 VGND.n334 121.493
R893 VGND.n213 VGND.t374 118.005
R894 VGND.n199 VGND.t339 118.005
R895 VGND.n461 VGND.t322 118.005
R896 VGND.n446 VGND.t331 118.005
R897 VGND.n690 VGND.t311 118.005
R898 VGND.n669 VGND.t313 118.005
R899 VGND.n776 VGND.t215 118.005
R900 VGND.n762 VGND.t260 118.005
R901 VGND.n974 VGND.t355 118.005
R902 VGND.n959 VGND.t367 118.005
R903 VGND.n911 VGND.t247 118.005
R904 VGND.n896 VGND.t232 118.005
R905 VGND.n287 VGND.t348 118.005
R906 VGND.n273 VGND.t341 118.005
R907 VGND.n406 VGND.t229 118.005
R908 VGND.n391 VGND.t281 118.005
R909 VGND.n249 VGND.n165 113.481
R910 VGND.n534 VGND.n78 113.481
R911 VGND.n819 VGND.n818 113.481
R912 VGND.n948 VGND.n947 113.481
R913 VGND.n1049 VGND.n1048 113.481
R914 VGND.n323 VGND.n139 113.481
R915 VGND.n380 VGND.n379 113.481
R916 VGND VGND.t24 111.335
R917 VGND.t137 VGND.t82 110.659
R918 VGND.t29 VGND.t137 110.659
R919 VGND.t80 VGND.t29 110.659
R920 VGND.t84 VGND.t80 110.659
R921 VGND.t26 VGND.t84 110.659
R922 VGND.t453 VGND 109.805
R923 VGND.t168 VGND.t164 108.898
R924 VGND.t164 VGND.t166 108.898
R925 VGND.t166 VGND.t451 108.898
R926 VGND.t451 VGND.t34 108.898
R927 VGND.t34 VGND.t45 108.898
R928 VGND.n259 VGND.n75 108.686
R929 VGND.n214 VGND.t300 104.028
R930 VGND.n212 VGND.t235 104.028
R931 VGND.n211 VGND.t270 104.028
R932 VGND.n197 VGND.t360 104.028
R933 VGND.n203 VGND.t304 104.028
R934 VGND.n198 VGND.t241 104.028
R935 VGND.n462 VGND.t352 104.028
R936 VGND.n460 VGND.t308 104.028
R937 VGND.n459 VGND.t297 104.028
R938 VGND.n444 VGND.t250 104.028
R939 VGND.n450 VGND.t357 104.028
R940 VGND.n445 VGND.t365 104.028
R941 VGND.n691 VGND.t206 104.028
R942 VGND.n689 VGND.t218 104.028
R943 VGND.n688 VGND.t362 104.028
R944 VGND.n667 VGND.t292 104.028
R945 VGND.n673 VGND.t212 104.028
R946 VGND.n668 VGND.t221 104.028
R947 VGND.n777 VGND.t253 104.028
R948 VGND.n775 VGND.t263 104.028
R949 VGND.n774 VGND.t376 104.028
R950 VGND.n760 VGND.t325 104.028
R951 VGND.n766 VGND.t278 104.028
R952 VGND.n761 VGND.t306 104.028
R953 VGND.n975 VGND.t266 104.028
R954 VGND.n973 VGND.t210 104.028
R955 VGND.n972 VGND.t238 104.028
R956 VGND.n957 VGND.t337 104.028
R957 VGND.n963 VGND.t275 104.028
R958 VGND.n958 VGND.t287 104.028
R959 VGND.n912 VGND.t334 104.028
R960 VGND.n910 VGND.t290 104.028
R961 VGND.n909 VGND.t226 104.028
R962 VGND.n894 VGND.t372 104.028
R963 VGND.n900 VGND.t345 104.028
R964 VGND.n895 VGND.t318 104.028
R965 VGND.n288 VGND.t256 104.028
R966 VGND.n286 VGND.t369 104.028
R967 VGND.n285 VGND.t328 104.028
R968 VGND.n271 VGND.t272 104.028
R969 VGND.n277 VGND.t284 104.028
R970 VGND.n272 VGND.t244 104.028
R971 VGND.n407 VGND.t315 104.028
R972 VGND.n405 VGND.t320 104.028
R973 VGND.n404 VGND.t295 104.028
R974 VGND.n389 VGND.t224 104.028
R975 VGND.n395 VGND.t343 104.028
R976 VGND.n390 VGND.t350 104.028
R977 VGND.n1026 VGND.n1025 101.547
R978 VGND.t0 VGND.t13 100.38
R979 VGND.t13 VGND.t9 100.38
R980 VGND.t9 VGND.t2 100.38
R981 VGND.t2 VGND.t16 100.38
R982 VGND.t16 VGND.t4 100.38
R983 VGND.t4 VGND.t7 100.38
R984 VGND.t7 VGND.t11 100.38
R985 VGND.t402 VGND.t404 100.38
R986 VGND.t404 VGND.t400 100.38
R987 VGND.n364 VGND.n363 99.7813
R988 VGND.t45 VGND.t449 99.3969
R989 VGND.t11 VGND.n262 97.9907
R990 VGND.t24 VGND.t135 95.4304
R991 VGND.t449 VGND.t453 94.1181
R992 VGND.n737 VGND.n727 93.189
R993 VGND.n357 VGND.n356 92.9264
R994 VGND.n1039 VGND.n58 92.9264
R995 VGND.n1035 VGND.n1034 92.9264
R996 VGND.n754 VGND.n721 92.9264
R997 VGND.n601 VGND.n595 92.9264
R998 VGND.n610 VGND.n603 92.9264
R999 VGND.n564 VGND.n563 92.9264
R1000 VGND.n1006 VGND.n556 92.9264
R1001 VGND.n733 VGND.n732 92.9264
R1002 VGND.n832 VGND.n568 92.9264
R1003 VGND.n575 VGND.n574 92.9264
R1004 VGND.n147 VGND.n146 92.9264
R1005 VGND.n520 VGND.n94 92.9264
R1006 VGND.n352 VGND.n351 92.9264
R1007 VGND.n1062 VGND.n29 92.9264
R1008 VGND.n375 VGND.n374 92.62
R1009 VGND.t135 VGND.t26 92.274
R1010 VGND.n543 VGND.t177 92.2476
R1011 VGND.n528 VGND.n527 92.0281
R1012 VGND.n746 VGND.n740 88.4348
R1013 VGND.n213 VGND.t375 87.6949
R1014 VGND.n461 VGND.t324 87.6949
R1015 VGND.n690 VGND.t312 87.6949
R1016 VGND.n776 VGND.t217 87.6949
R1017 VGND.n974 VGND.t356 87.6949
R1018 VGND.n911 VGND.t249 87.6949
R1019 VGND.n287 VGND.t349 87.6949
R1020 VGND.n406 VGND.t231 87.6949
R1021 VGND.n199 VGND.t340 87.5315
R1022 VGND.n446 VGND.t333 87.5315
R1023 VGND.n669 VGND.t314 87.5315
R1024 VGND.n762 VGND.t262 87.5315
R1025 VGND.n959 VGND.t368 87.5315
R1026 VGND.n896 VGND.t234 87.5315
R1027 VGND.n273 VGND.t342 87.5315
R1028 VGND.n391 VGND.t283 87.5315
R1029 VGND.n363 VGND.n334 82.4308
R1030 VGND.n256 VGND.n255 80.224
R1031 VGND.n531 VGND.n530 80.224
R1032 VGND.n823 VGND.n822 80.224
R1033 VGND.n1053 VGND.n1052 80.224
R1034 VGND.n330 VGND.n329 80.224
R1035 VGND.n372 VGND.n371 80.224
R1036 VGND.t177 VGND 79.8654
R1037 VGND.t28 VGND.n334 78.5719
R1038 VGND.t72 VGND.n225 77.0353
R1039 VGND.t51 VGND.n443 77.0353
R1040 VGND.t193 VGND.n686 77.0353
R1041 VGND.t194 VGND.n788 77.0353
R1042 VGND.t152 VGND.n956 77.0353
R1043 VGND.t195 VGND.n893 77.0353
R1044 VGND.t448 VGND.n299 77.0353
R1045 VGND.t382 VGND.n388 77.0353
R1046 VGND.n163 VGND.n162 67.8728
R1047 VGND.n84 VGND.n81 67.8728
R1048 VGND.n821 VGND.n594 67.8728
R1049 VGND.n945 VGND.n944 67.8728
R1050 VGND.n1051 VGND.n40 67.8728
R1051 VGND.n137 VGND.n136 67.8728
R1052 VGND.n366 VGND.n122 67.8728
R1053 VGND.n132 VGND.n34 65.486
R1054 VGND.n52 VGND.n51 65.486
R1055 VGND.n590 VGND.n589 65.486
R1056 VGND.n85 VGND.n75 65.486
R1057 VGND.n158 VGND.n64 65.486
R1058 VGND.n1019 VGND.n540 65.486
R1059 VGND.n1033 VGND.n1032 65.0005
R1060 VGND.n62 VGND.n57 65.0005
R1061 VGND.n751 VGND.n723 65.0005
R1062 VGND.n599 VGND.n598 65.0005
R1063 VGND.n608 VGND.n607 65.0005
R1064 VGND.n562 VGND.n561 65.0005
R1065 VGND.n555 VGND.n554 65.0005
R1066 VGND.n731 VGND.n730 65.0005
R1067 VGND.n829 VGND.n570 65.0005
R1068 VGND.n746 VGND.n745 65.0005
R1069 VGND.n745 VGND.n744 65.0005
R1070 VGND.n573 VGND.n572 65.0005
R1071 VGND.n145 VGND.n144 65.0005
R1072 VGND.n151 VGND.n93 65.0005
R1073 VGND.n350 VGND.n349 65.0005
R1074 VGND.n341 VGND.n338 65.0005
R1075 VGND.n1059 VGND.n31 65.0005
R1076 VGND.n260 VGND.n259 64.2492
R1077 VGND VGND.t55 64.1195
R1078 VGND.n1034 VGND.n1033 59.3637
R1079 VGND.n58 VGND.n57 59.3637
R1080 VGND.n723 VGND.n721 59.3637
R1081 VGND.n599 VGND.n595 59.3637
R1082 VGND.n608 VGND.n603 59.3637
R1083 VGND.n563 VGND.n562 59.3637
R1084 VGND.n556 VGND.n555 59.3637
R1085 VGND.n732 VGND.n731 59.3637
R1086 VGND.n570 VGND.n568 59.3637
R1087 VGND.n574 VGND.n573 59.3637
R1088 VGND.n147 VGND.n145 59.3637
R1089 VGND.n94 VGND.n93 59.3637
R1090 VGND.n351 VGND.n350 59.3637
R1091 VGND.n357 VGND.n338 59.3637
R1092 VGND.n31 VGND.n29 59.3637
R1093 VGND.n346 VGND.t127 58.4716
R1094 VGND.t430 VGND.n525 57.983
R1095 VGND.t57 VGND.t53 54.9596
R1096 VGND.t141 VGND.t57 54.9596
R1097 VGND.t143 VGND.t141 54.9596
R1098 VGND.n361 VGND.t143 48.4169
R1099 VGND.n362 VGND 43.8369
R1100 VGND.n618 VGND 42.3499
R1101 VGND.n865 VGND 42.3499
R1102 VGND.n220 VGND.t145 41.4291
R1103 VGND.n220 VGND.t271 41.4291
R1104 VGND.t237 VGND.n217 41.4291
R1105 VGND.n217 VGND.t302 41.4291
R1106 VGND.t271 VGND.n219 41.4291
R1107 VGND.n219 VGND.t237 41.4291
R1108 VGND.n222 VGND.t151 41.4291
R1109 VGND.n222 VGND.t150 41.4291
R1110 VGND.n206 VGND.t361 41.4291
R1111 VGND.n206 VGND.t147 41.4291
R1112 VGND.n205 VGND.t305 41.4291
R1113 VGND.t361 VGND.n205 41.4291
R1114 VGND.n201 VGND.t243 41.4291
R1115 VGND.n201 VGND.t305 41.4291
R1116 VGND.n208 VGND.t149 41.4291
R1117 VGND.n208 VGND.t148 41.4291
R1118 VGND.n468 VGND.t98 41.4291
R1119 VGND.n468 VGND.t299 41.4291
R1120 VGND.t310 VGND.n465 41.4291
R1121 VGND.n465 VGND.t353 41.4291
R1122 VGND.t299 VGND.n467 41.4291
R1123 VGND.n467 VGND.t310 41.4291
R1124 VGND.n470 VGND.t108 41.4291
R1125 VGND.n470 VGND.t100 41.4291
R1126 VGND.n453 VGND.t252 41.4291
R1127 VGND.n453 VGND.t102 41.4291
R1128 VGND.n452 VGND.t359 41.4291
R1129 VGND.t252 VGND.n452 41.4291
R1130 VGND.n448 VGND.t366 41.4291
R1131 VGND.n448 VGND.t359 41.4291
R1132 VGND.n455 VGND.t104 41.4291
R1133 VGND.n455 VGND.t106 41.4291
R1134 VGND.n697 VGND.t416 41.4291
R1135 VGND.n697 VGND.t364 41.4291
R1136 VGND.t220 VGND.n694 41.4291
R1137 VGND.n694 VGND.t208 41.4291
R1138 VGND.t364 VGND.n696 41.4291
R1139 VGND.n696 VGND.t220 41.4291
R1140 VGND.n699 VGND.t410 41.4291
R1141 VGND.n699 VGND.t414 41.4291
R1142 VGND.n676 VGND.t294 41.4291
R1143 VGND.n676 VGND.t417 41.4291
R1144 VGND.n675 VGND.t214 41.4291
R1145 VGND.t294 VGND.n675 41.4291
R1146 VGND.n671 VGND.t223 41.4291
R1147 VGND.n671 VGND.t214 41.4291
R1148 VGND.n678 VGND.t419 41.4291
R1149 VGND.n678 VGND.t412 41.4291
R1150 VGND.n783 VGND.t445 41.4291
R1151 VGND.n783 VGND.t378 41.4291
R1152 VGND.t265 VGND.n780 41.4291
R1153 VGND.n780 VGND.t254 41.4291
R1154 VGND.t378 VGND.n782 41.4291
R1155 VGND.n782 VGND.t265 41.4291
R1156 VGND.n785 VGND.t441 41.4291
R1157 VGND.n785 VGND.t444 41.4291
R1158 VGND.n769 VGND.t327 41.4291
R1159 VGND.n769 VGND.t447 41.4291
R1160 VGND.n768 VGND.t280 41.4291
R1161 VGND.t327 VGND.n768 41.4291
R1162 VGND.n764 VGND.t307 41.4291
R1163 VGND.n764 VGND.t280 41.4291
R1164 VGND.n771 VGND.t439 41.4291
R1165 VGND.n771 VGND.t442 41.4291
R1166 VGND.n981 VGND.t467 41.4291
R1167 VGND.n981 VGND.t240 41.4291
R1168 VGND.t211 VGND.n978 41.4291
R1169 VGND.n978 VGND.t268 41.4291
R1170 VGND.t240 VGND.n980 41.4291
R1171 VGND.n980 VGND.t211 41.4291
R1172 VGND.n983 VGND.t465 41.4291
R1173 VGND.n983 VGND.t466 41.4291
R1174 VGND.n966 VGND.t338 41.4291
R1175 VGND.n966 VGND.t468 41.4291
R1176 VGND.n965 VGND.t277 41.4291
R1177 VGND.t338 VGND.n965 41.4291
R1178 VGND.n961 VGND.t289 41.4291
R1179 VGND.n961 VGND.t277 41.4291
R1180 VGND.n968 VGND.t464 41.4291
R1181 VGND.n968 VGND.t463 41.4291
R1182 VGND.n918 VGND.t155 41.4291
R1183 VGND.n918 VGND.t228 41.4291
R1184 VGND.t291 VGND.n915 41.4291
R1185 VGND.n915 VGND.t335 41.4291
R1186 VGND.t228 VGND.n917 41.4291
R1187 VGND.n917 VGND.t291 41.4291
R1188 VGND.n920 VGND.t161 41.4291
R1189 VGND.n920 VGND.t162 41.4291
R1190 VGND.n903 VGND.t373 41.4291
R1191 VGND.n903 VGND.t156 41.4291
R1192 VGND.n902 VGND.t347 41.4291
R1193 VGND.t373 VGND.n902 41.4291
R1194 VGND.n898 VGND.t319 41.4291
R1195 VGND.n898 VGND.t347 41.4291
R1196 VGND.n905 VGND.t160 41.4291
R1197 VGND.n905 VGND.t158 41.4291
R1198 VGND.n294 VGND.t189 41.4291
R1199 VGND.n294 VGND.t330 41.4291
R1200 VGND.t371 VGND.n291 41.4291
R1201 VGND.n291 VGND.t258 41.4291
R1202 VGND.t330 VGND.n293 41.4291
R1203 VGND.n293 VGND.t371 41.4291
R1204 VGND.n296 VGND.t187 41.4291
R1205 VGND.n296 VGND.t185 41.4291
R1206 VGND.n280 VGND.t274 41.4291
R1207 VGND.n280 VGND.t191 41.4291
R1208 VGND.n279 VGND.t286 41.4291
R1209 VGND.t274 VGND.n279 41.4291
R1210 VGND.n275 VGND.t246 41.4291
R1211 VGND.n275 VGND.t286 41.4291
R1212 VGND.n282 VGND.t183 41.4291
R1213 VGND.n282 VGND.t181 41.4291
R1214 VGND.n413 VGND.t398 41.4291
R1215 VGND.n413 VGND.t296 41.4291
R1216 VGND.t321 VGND.n410 41.4291
R1217 VGND.n410 VGND.t316 41.4291
R1218 VGND.t296 VGND.n412 41.4291
R1219 VGND.n412 VGND.t321 41.4291
R1220 VGND.n415 VGND.t396 41.4291
R1221 VGND.n415 VGND.t399 41.4291
R1222 VGND.n398 VGND.t225 41.4291
R1223 VGND.n398 VGND.t394 41.4291
R1224 VGND.n397 VGND.t344 41.4291
R1225 VGND.t225 VGND.n397 41.4291
R1226 VGND.n393 VGND.t351 41.4291
R1227 VGND.n393 VGND.t344 41.4291
R1228 VGND.n400 VGND.t395 41.4291
R1229 VGND.n400 VGND.t397 41.4291
R1230 VGND.t172 VGND.n542 37.7835
R1231 VGND.t53 VGND.n360 36.6399
R1232 VGND.n250 VGND.n249 36.4805
R1233 VGND.n79 VGND.n78 36.4805
R1234 VGND.n819 VGND.n811 36.4805
R1235 VGND.n948 VGND.n946 36.4805
R1236 VGND.n1049 VGND.n42 36.4805
R1237 VGND.n324 VGND.n323 36.4805
R1238 VGND.n380 VGND.n123 36.4805
R1239 VGND VGND.n171 35.197
R1240 VGND VGND.n99 35.197
R1241 VGND VGND.n644 35.197
R1242 VGND VGND.n838 35.197
R1243 VGND VGND.n494 35.197
R1244 VGND VGND.n5 35.197
R1245 VGND.n175 VGND.n174 34.6358
R1246 VGND.n188 VGND.n187 34.6358
R1247 VGND.n184 VGND.n183 34.6358
R1248 VGND.n103 VGND.n102 34.6358
R1249 VGND.n116 VGND.n115 34.6358
R1250 VGND.n112 VGND.n111 34.6358
R1251 VGND.n622 VGND.n621 34.6358
R1252 VGND.n635 VGND.n634 34.6358
R1253 VGND.n631 VGND.n630 34.6358
R1254 VGND.n648 VGND.n647 34.6358
R1255 VGND.n661 VGND.n660 34.6358
R1256 VGND.n657 VGND.n656 34.6358
R1257 VGND.n869 VGND.n868 34.6358
R1258 VGND.n882 VGND.n881 34.6358
R1259 VGND.n878 VGND.n877 34.6358
R1260 VGND.n842 VGND.n841 34.6358
R1261 VGND.n855 VGND.n854 34.6358
R1262 VGND.n851 VGND.n850 34.6358
R1263 VGND.n498 VGND.n497 34.6358
R1264 VGND.n511 VGND.n510 34.6358
R1265 VGND.n507 VGND.n506 34.6358
R1266 VGND.n9 VGND.n8 34.6358
R1267 VGND.n22 VGND.n21 34.6358
R1268 VGND.n18 VGND.n17 34.6358
R1269 VGND.n360 VGND.t400 33.4606
R1270 VGND.n190 VGND.n189 32.0005
R1271 VGND.n118 VGND.n117 32.0005
R1272 VGND.n637 VGND.n636 32.0005
R1273 VGND.n663 VGND.n662 32.0005
R1274 VGND.n884 VGND.n883 32.0005
R1275 VGND.n857 VGND.n856 32.0005
R1276 VGND.n513 VGND.n512 32.0005
R1277 VGND.n24 VGND.n23 32.0005
R1278 VGND.n826 VGND.n52 31.5543
R1279 VGND.n190 VGND.n176 31.2476
R1280 VGND.n118 VGND.n104 31.2476
R1281 VGND.n637 VGND.n623 31.2476
R1282 VGND.n663 VGND.n649 31.2476
R1283 VGND.n884 VGND.n870 31.2476
R1284 VGND.n857 VGND.n843 31.2476
R1285 VGND.n513 VGND.n499 31.2476
R1286 VGND.n24 VGND.n10 31.2476
R1287 VGND.n621 VGND.n617 30.1181
R1288 VGND.n868 VGND.n864 30.1181
R1289 VGND.t110 VGND 28.0716
R1290 VGND VGND.t66 27.836
R1291 VGND.n245 VGND.n244 26.2219
R1292 VGND.n473 VGND.n472 26.2219
R1293 VGND.n702 VGND.n701 26.2219
R1294 VGND.n808 VGND.n807 26.2219
R1295 VGND.n986 VGND.n985 26.2219
R1296 VGND.n923 VGND.n922 26.2219
R1297 VGND.n319 VGND.n318 26.2219
R1298 VGND.n418 VGND.n417 26.2219
R1299 VGND.n187 VGND.n179 25.977
R1300 VGND.n115 VGND.n107 25.977
R1301 VGND.n634 VGND.n626 25.977
R1302 VGND.n660 VGND.n652 25.977
R1303 VGND.n881 VGND.n873 25.977
R1304 VGND.n854 VGND.n846 25.977
R1305 VGND.n510 VGND.n502 25.977
R1306 VGND.n21 VGND.n13 25.977
R1307 VGND.n265 VGND.n264 25.0956
R1308 VGND.n170 VGND.t14 24.9236
R1309 VGND.n170 VGND.t10 24.9236
R1310 VGND.n177 VGND.t3 24.9236
R1311 VGND.n177 VGND.t17 24.9236
R1312 VGND.n178 VGND.t5 24.9236
R1313 VGND.n178 VGND.t8 24.9236
R1314 VGND.n98 VGND.t134 24.9236
R1315 VGND.n98 VGND.t115 24.9236
R1316 VGND.n105 VGND.t117 24.9236
R1317 VGND.n105 VGND.t132 24.9236
R1318 VGND.n106 VGND.t113 24.9236
R1319 VGND.n106 VGND.t130 24.9236
R1320 VGND.n616 VGND.t176 24.9236
R1321 VGND.n616 VGND.t121 24.9236
R1322 VGND.n624 VGND.t126 24.9236
R1323 VGND.n624 VGND.t71 24.9236
R1324 VGND.n625 VGND.t124 24.9236
R1325 VGND.n625 VGND.t173 24.9236
R1326 VGND.n643 VGND.t462 24.9236
R1327 VGND.n643 VGND.t22 24.9236
R1328 VGND.n650 VGND.t423 24.9236
R1329 VGND.n650 VGND.t460 24.9236
R1330 VGND.n651 VGND.t20 24.9236
R1331 VGND.n651 VGND.t475 24.9236
R1332 VGND.n863 VGND.t138 24.9236
R1333 VGND.n863 VGND.t30 24.9236
R1334 VGND.n871 VGND.t81 24.9236
R1335 VGND.n871 VGND.t85 24.9236
R1336 VGND.n872 VGND.t27 24.9236
R1337 VGND.n872 VGND.t136 24.9236
R1338 VGND.n837 VGND.t165 24.9236
R1339 VGND.n837 VGND.t167 24.9236
R1340 VGND.n844 VGND.t452 24.9236
R1341 VGND.n844 VGND.t35 24.9236
R1342 VGND.n845 VGND.t46 24.9236
R1343 VGND.n845 VGND.t450 24.9236
R1344 VGND.n493 VGND.t435 24.9236
R1345 VGND.n493 VGND.t48 24.9236
R1346 VGND.n500 VGND.t50 24.9236
R1347 VGND.n500 VGND.t437 24.9236
R1348 VGND.n501 VGND.t429 24.9236
R1349 VGND.n501 VGND.t433 24.9236
R1350 VGND.n4 VGND.t405 24.9236
R1351 VGND.n4 VGND.t401 24.9236
R1352 VGND.n11 VGND.t54 24.9236
R1353 VGND.n11 VGND.t58 24.9236
R1354 VGND.n12 VGND.t142 24.9236
R1355 VGND.n12 VGND.t144 24.9236
R1356 VGND.t127 VGND.t133 24.0614
R1357 VGND.t133 VGND.t114 24.0614
R1358 VGND.t114 VGND.t116 24.0614
R1359 VGND.t116 VGND.t131 24.0614
R1360 VGND.t131 VGND.t112 24.0614
R1361 VGND.t112 VGND.t129 24.0614
R1362 VGND.t129 VGND.t110 24.0614
R1363 VGND.n1022 VGND.n70 23.993
R1364 VGND.t434 VGND.t430 23.8595
R1365 VGND.t47 VGND.t434 23.8595
R1366 VGND.t49 VGND.t47 23.8595
R1367 VGND.t436 VGND.t49 23.8595
R1368 VGND.t428 VGND.t436 23.8595
R1369 VGND.t432 VGND.t428 23.8595
R1370 VGND.t66 VGND.t432 23.8595
R1371 VGND.n826 VGND.n583 23.8559
R1372 VGND.n378 VGND.n377 23.4005
R1373 VGND.n377 VGND.t389 23.4005
R1374 VGND.n376 VGND.n123 23.4005
R1375 VGND.t389 VGND.n376 23.4005
R1376 VGND.n327 VGND.n326 23.4005
R1377 VGND.n326 VGND.t469 23.4005
R1378 VGND.n325 VGND.n324 23.4005
R1379 VGND.t469 VGND.n325 23.4005
R1380 VGND.n47 VGND.n43 23.4005
R1381 VGND.t62 VGND.n47 23.4005
R1382 VGND.n44 VGND.n42 23.4005
R1383 VGND.t62 VGND.n44 23.4005
R1384 VGND.n816 VGND.n812 23.4005
R1385 VGND.n816 VGND.t386 23.4005
R1386 VGND.n813 VGND.n811 23.4005
R1387 VGND.t386 VGND.n813 23.4005
R1388 VGND.n253 VGND.n252 23.4005
R1389 VGND.n252 VGND.t88 23.4005
R1390 VGND.n251 VGND.n250 23.4005
R1391 VGND.t88 VGND.n251 23.4005
R1392 VGND.n1022 VGND.t59 23.4005
R1393 VGND.n946 VGND.n72 23.4005
R1394 VGND.t59 VGND.n72 23.4005
R1395 VGND.n533 VGND.n77 23.4005
R1396 VGND.n77 VGND.t383 23.4005
R1397 VGND.n79 VGND.n76 23.4005
R1398 VGND.n76 VGND.t383 23.4005
R1399 VGND.n630 VGND.n629 23.3417
R1400 VGND.n877 VGND.n876 23.3417
R1401 VGND.n1011 VGND.n1010 22.6809
R1402 VGND.n132 VGND.n129 21.6084
R1403 VGND.n51 VGND.n36 21.6084
R1404 VGND.n590 VGND.n585 21.6084
R1405 VGND.n85 VGND.n83 21.6084
R1406 VGND.n158 VGND.n155 21.6084
R1407 VGND.n540 VGND.n67 21.6084
R1408 VGND.n227 VGND.n225 20.8934
R1409 VGND.n234 VGND.n224 20.8934
R1410 VGND.n478 VGND.n443 20.8934
R1411 VGND.n475 VGND.n442 20.8934
R1412 VGND.n707 VGND.n686 20.8934
R1413 VGND.n704 VGND.n685 20.8934
R1414 VGND.n790 VGND.n788 20.8934
R1415 VGND.n797 VGND.n787 20.8934
R1416 VGND.n991 VGND.n956 20.8934
R1417 VGND.n988 VGND.n955 20.8934
R1418 VGND.n928 VGND.n893 20.8934
R1419 VGND.n925 VGND.n892 20.8934
R1420 VGND.n301 VGND.n299 20.8934
R1421 VGND.n308 VGND.n298 20.8934
R1422 VGND.n423 VGND.n388 20.8934
R1423 VGND.n420 VGND.n387 20.8934
R1424 VGND.n629 VGND.n628 20.5946
R1425 VGND.n876 VGND.n875 20.5946
R1426 VGND.n262 VGND 19.1205
R1427 VGND.n174 VGND.n171 18.824
R1428 VGND.n102 VGND.n99 18.824
R1429 VGND.n647 VGND.n644 18.824
R1430 VGND.n841 VGND.n838 18.824
R1431 VGND.n497 VGND.n494 18.824
R1432 VGND.n8 VGND.n5 18.824
R1433 VGND.n374 VGND.n334 14.2936
R1434 VGND.n366 VGND.n365 13.6052
R1435 VGND.n370 VGND.n364 13.6052
R1436 VGND.n136 VGND.n130 13.6052
R1437 VGND.n131 VGND.n129 13.6052
R1438 VGND.n40 VGND.n37 13.6052
R1439 VGND.n38 VGND.n36 13.6052
R1440 VGND.n594 VGND.n586 13.6052
R1441 VGND.n587 VGND.n585 13.6052
R1442 VGND.n89 VGND.n84 13.6052
R1443 VGND.n83 VGND.n82 13.6052
R1444 VGND.n162 VGND.n156 13.6052
R1445 VGND.n157 VGND.n155 13.6052
R1446 VGND.n944 VGND.n68 13.6052
R1447 VGND.n69 VGND.n67 13.6052
R1448 VGND.n183 VGND.n182 13.5534
R1449 VGND.n111 VGND.n110 13.5534
R1450 VGND.n656 VGND.n655 13.5534
R1451 VGND.n850 VGND.n849 13.5534
R1452 VGND.n506 VGND.n505 13.5534
R1453 VGND.n17 VGND.n16 13.5534
R1454 VGND.n254 VGND.n164 13.177
R1455 VGND.n532 VGND.n80 13.177
R1456 VGND.n814 VGND.n588 13.177
R1457 VGND.n45 VGND.n39 13.177
R1458 VGND.n328 VGND.n138 13.177
R1459 VGND.n126 VGND.n125 13.177
R1460 VGND.n356 VGND 11.4981
R1461 VGND.n1039 VGND 11.4981
R1462 VGND VGND.n1035 11.4981
R1463 VGND VGND.n754 11.4981
R1464 VGND VGND.n601 11.4981
R1465 VGND VGND.n610 11.4981
R1466 VGND VGND.n564 11.4981
R1467 VGND.n1006 VGND 11.4981
R1468 VGND.n733 VGND 11.4981
R1469 VGND VGND.n832 11.4981
R1470 VGND.n740 VGND 11.4981
R1471 VGND.n575 VGND 11.4981
R1472 VGND.n146 VGND 11.4981
R1473 VGND.n520 VGND 11.4981
R1474 VGND VGND.n352 11.4981
R1475 VGND VGND.n1062 11.4981
R1476 VGND.n182 VGND.n181 11.1829
R1477 VGND.n110 VGND.n109 11.1829
R1478 VGND.n655 VGND.n654 11.1829
R1479 VGND.n849 VGND.n848 11.1829
R1480 VGND.n505 VGND.n504 11.1829
R1481 VGND.n16 VGND.n15 11.1829
R1482 VGND.n1044 VGND.n1043 11.1086
R1483 VGND.n1025 VGND.n1024 10.2529
R1484 VGND.n172 VGND.n171 9.3005
R1485 VGND.n174 VGND.n173 9.3005
R1486 VGND.n175 VGND.n168 9.3005
R1487 VGND.n191 VGND.n190 9.3005
R1488 VGND.n188 VGND.n169 9.3005
R1489 VGND.n187 VGND.n186 9.3005
R1490 VGND.n185 VGND.n184 9.3005
R1491 VGND.n183 VGND.n180 9.3005
R1492 VGND.n100 VGND.n99 9.3005
R1493 VGND.n102 VGND.n101 9.3005
R1494 VGND.n103 VGND.n96 9.3005
R1495 VGND.n119 VGND.n118 9.3005
R1496 VGND.n116 VGND.n97 9.3005
R1497 VGND.n115 VGND.n114 9.3005
R1498 VGND.n113 VGND.n112 9.3005
R1499 VGND.n111 VGND.n108 9.3005
R1500 VGND.n619 VGND.n618 9.3005
R1501 VGND.n621 VGND.n620 9.3005
R1502 VGND.n622 VGND.n614 9.3005
R1503 VGND.n638 VGND.n637 9.3005
R1504 VGND.n635 VGND.n615 9.3005
R1505 VGND.n634 VGND.n633 9.3005
R1506 VGND.n632 VGND.n631 9.3005
R1507 VGND.n630 VGND.n627 9.3005
R1508 VGND.n645 VGND.n644 9.3005
R1509 VGND.n647 VGND.n646 9.3005
R1510 VGND.n648 VGND.n641 9.3005
R1511 VGND.n664 VGND.n663 9.3005
R1512 VGND.n661 VGND.n642 9.3005
R1513 VGND.n660 VGND.n659 9.3005
R1514 VGND.n658 VGND.n657 9.3005
R1515 VGND.n656 VGND.n653 9.3005
R1516 VGND.n866 VGND.n865 9.3005
R1517 VGND.n868 VGND.n867 9.3005
R1518 VGND.n869 VGND.n861 9.3005
R1519 VGND.n885 VGND.n884 9.3005
R1520 VGND.n882 VGND.n862 9.3005
R1521 VGND.n881 VGND.n880 9.3005
R1522 VGND.n879 VGND.n878 9.3005
R1523 VGND.n877 VGND.n874 9.3005
R1524 VGND.n839 VGND.n838 9.3005
R1525 VGND.n841 VGND.n840 9.3005
R1526 VGND.n842 VGND.n835 9.3005
R1527 VGND.n858 VGND.n857 9.3005
R1528 VGND.n855 VGND.n836 9.3005
R1529 VGND.n854 VGND.n853 9.3005
R1530 VGND.n852 VGND.n851 9.3005
R1531 VGND.n850 VGND.n847 9.3005
R1532 VGND.n495 VGND.n494 9.3005
R1533 VGND.n497 VGND.n496 9.3005
R1534 VGND.n498 VGND.n491 9.3005
R1535 VGND.n514 VGND.n513 9.3005
R1536 VGND.n511 VGND.n492 9.3005
R1537 VGND.n510 VGND.n509 9.3005
R1538 VGND.n508 VGND.n507 9.3005
R1539 VGND.n506 VGND.n503 9.3005
R1540 VGND.n6 VGND.n5 9.3005
R1541 VGND.n8 VGND.n7 9.3005
R1542 VGND.n9 VGND.n2 9.3005
R1543 VGND.n25 VGND.n24 9.3005
R1544 VGND.n22 VGND.n3 9.3005
R1545 VGND.n21 VGND.n20 9.3005
R1546 VGND.n19 VGND.n18 9.3005
R1547 VGND.n17 VGND.n14 9.3005
R1548 VGND.n184 VGND.n179 8.65932
R1549 VGND.n112 VGND.n107 8.65932
R1550 VGND.n631 VGND.n626 8.65932
R1551 VGND.n657 VGND.n652 8.65932
R1552 VGND.n878 VGND.n873 8.65932
R1553 VGND.n851 VGND.n846 8.65932
R1554 VGND.n507 VGND.n502 8.65932
R1555 VGND.n18 VGND.n13 8.65932
R1556 VGND.n726 VGND.n724 8.57205
R1557 VGND.n232 VGND.n231 8.23994
R1558 VGND.n231 VGND.n230 8.23994
R1559 VGND.n242 VGND.n241 8.23994
R1560 VGND.n243 VGND.n242 8.23994
R1561 VGND.n480 VGND.n479 8.23994
R1562 VGND.n481 VGND.n480 8.23994
R1563 VGND.n484 VGND.n483 8.23994
R1564 VGND.n483 VGND.n482 8.23994
R1565 VGND.n709 VGND.n708 8.23994
R1566 VGND.n710 VGND.n709 8.23994
R1567 VGND.n713 VGND.n712 8.23994
R1568 VGND.n712 VGND.n711 8.23994
R1569 VGND.n795 VGND.n794 8.23994
R1570 VGND.n794 VGND.n793 8.23994
R1571 VGND.n805 VGND.n804 8.23994
R1572 VGND.n806 VGND.n805 8.23994
R1573 VGND.n993 VGND.n992 8.23994
R1574 VGND.n994 VGND.n993 8.23994
R1575 VGND.n997 VGND.n996 8.23994
R1576 VGND.n996 VGND.n995 8.23994
R1577 VGND.n930 VGND.n929 8.23994
R1578 VGND.n931 VGND.n930 8.23994
R1579 VGND.n934 VGND.n933 8.23994
R1580 VGND.n933 VGND.n932 8.23994
R1581 VGND.n306 VGND.n305 8.23994
R1582 VGND.n305 VGND.n304 8.23994
R1583 VGND.n316 VGND.n315 8.23994
R1584 VGND.n317 VGND.n316 8.23994
R1585 VGND.n425 VGND.n424 8.23994
R1586 VGND.n426 VGND.n425 8.23994
R1587 VGND.n429 VGND.n428 8.23994
R1588 VGND.n428 VGND.n427 8.23994
R1589 VGND.n1024 VGND.n71 7.76749
R1590 VGND.t55 VGND.n361 6.54325
R1591 VGND.n133 VGND.t438 6.2726
R1592 VGND.t153 VGND.n50 6.2726
R1593 VGND.n591 VGND.t39 6.2726
R1594 VGND.n88 VGND.t23 6.2726
R1595 VGND.n159 VGND.t192 6.2726
R1596 VGND.n941 VGND.t179 6.2726
R1597 VGND.n367 VGND.t28 5.66771
R1598 VGND.n757 VGND 5.54759
R1599 VGND.n566 VGND 4.6065
R1600 VGND.n618 VGND.n617 4.51815
R1601 VGND.n865 VGND.n864 4.51815
R1602 VGND.n255 VGND.n254 4.3205
R1603 VGND.n532 VGND.n531 4.3205
R1604 VGND.n822 VGND.n588 4.3205
R1605 VGND.n1052 VGND.n39 4.3205
R1606 VGND.n329 VGND.n328 4.3205
R1607 VGND.n371 VGND.n125 4.3205
R1608 VGND.n1066 VGND 3.54117
R1609 VGND.n756 VGND.n720 3.45067
R1610 VGND.n355 VGND.n354 3.45067
R1611 VGND.n1038 VGND.n1037 3.45067
R1612 VGND.n612 VGND.n602 3.45067
R1613 VGND.n1004 VGND.n565 3.45067
R1614 VGND.n834 VGND.n567 3.45067
R1615 VGND.n518 VGND.n95 3.45067
R1616 VGND.n1064 VGND.n28 3.45067
R1617 VGND.n176 VGND.n175 3.38874
R1618 VGND.n104 VGND.n103 3.38874
R1619 VGND.n623 VGND.n622 3.38874
R1620 VGND.n649 VGND.n648 3.38874
R1621 VGND.n870 VGND.n869 3.38874
R1622 VGND.n843 VGND.n842 3.38874
R1623 VGND.n499 VGND.n498 3.38874
R1624 VGND.n10 VGND.n9 3.38874
R1625 VGND.n1037 VGND.n1036 2.87883
R1626 VGND.n756 VGND.n755 2.87883
R1627 VGND.n612 VGND.n611 2.87883
R1628 VGND.n1005 VGND.n1004 2.87883
R1629 VGND.n834 VGND.n833 2.87883
R1630 VGND.n519 VGND.n518 2.87883
R1631 VGND.n354 VGND.n353 2.87883
R1632 VGND.n1064 VGND.n1063 2.87883
R1633 VGND.n189 VGND.n188 2.63579
R1634 VGND.n117 VGND.n116 2.63579
R1635 VGND.n636 VGND.n635 2.63579
R1636 VGND.n662 VGND.n661 2.63579
R1637 VGND.n883 VGND.n882 2.63579
R1638 VGND.n856 VGND.n855 2.63579
R1639 VGND.n512 VGND.n511 2.63579
R1640 VGND.n23 VGND.n22 2.63579
R1641 VGND.n1067 VGND 2.47583
R1642 VGND.n248 VGND.n163 2.45057
R1643 VGND.n436 VGND.n81 2.45057
R1644 VGND.n821 VGND.n820 2.45057
R1645 VGND.n949 VGND.n945 2.45057
R1646 VGND.n1051 VGND.n1050 2.45057
R1647 VGND.n322 VGND.n137 2.45057
R1648 VGND.n381 VGND.n122 2.45057
R1649 VGND.n1069 VGND 2.2565
R1650 VGND.n239 VGND.n228 2.09737
R1651 VGND.n239 VGND.n238 2.09737
R1652 VGND.n476 VGND.n439 2.09737
R1653 VGND.n486 VGND.n439 2.09737
R1654 VGND.n705 VGND.n682 2.09737
R1655 VGND.n715 VGND.n682 2.09737
R1656 VGND.n802 VGND.n791 2.09737
R1657 VGND.n802 VGND.n801 2.09737
R1658 VGND.n989 VGND.n952 2.09737
R1659 VGND.n999 VGND.n952 2.09737
R1660 VGND.n926 VGND.n889 2.09737
R1661 VGND.n936 VGND.n889 2.09737
R1662 VGND.n313 VGND.n302 2.09737
R1663 VGND.n313 VGND.n312 2.09737
R1664 VGND.n421 VGND.n384 2.09737
R1665 VGND.n431 VGND.n384 2.09737
R1666 VGND.n236 VGND.n228 2.09113
R1667 VGND.n476 VGND.n438 2.09113
R1668 VGND.n705 VGND.n681 2.09113
R1669 VGND.n799 VGND.n791 2.09113
R1670 VGND.n989 VGND.n951 2.09113
R1671 VGND.n926 VGND.n888 2.09113
R1672 VGND.n310 VGND.n302 2.09113
R1673 VGND.n421 VGND.n383 2.09113
R1674 VGND.n233 VGND.n232 1.93989
R1675 VGND.n479 VGND.n477 1.93989
R1676 VGND.n708 VGND.n706 1.93989
R1677 VGND.n796 VGND.n795 1.93989
R1678 VGND.n992 VGND.n990 1.93989
R1679 VGND.n929 VGND.n927 1.93989
R1680 VGND.n307 VGND.n306 1.93989
R1681 VGND.n424 VGND.n422 1.93989
R1682 VGND.n237 VGND.n236 1.72862
R1683 VGND.n487 VGND.n438 1.72862
R1684 VGND.n716 VGND.n681 1.72862
R1685 VGND.n800 VGND.n799 1.72862
R1686 VGND.n1000 VGND.n951 1.72862
R1687 VGND.n937 VGND.n888 1.72862
R1688 VGND.n311 VGND.n310 1.72862
R1689 VGND.n432 VGND.n383 1.72862
R1690 VGND.n193 VGND.n192 1.24162
R1691 VGND.n121 VGND.n120 1.24162
R1692 VGND.n640 VGND.n639 1.24162
R1693 VGND.n666 VGND.n665 1.24162
R1694 VGND.n887 VGND.n886 1.24162
R1695 VGND.n860 VGND.n859 1.24162
R1696 VGND.n516 VGND.n515 1.24162
R1697 VGND.n27 VGND.n26 1.24162
R1698 VGND.n724 VGND.t424 1.00615
R1699 VGND.n240 VGND.n227 0.970197
R1700 VGND.n241 VGND.n226 0.970197
R1701 VGND.n235 VGND.n234 0.970197
R1702 VGND.n478 VGND.n441 0.970197
R1703 VGND.n485 VGND.n484 0.970197
R1704 VGND.n475 VGND.n440 0.970197
R1705 VGND.n707 VGND.n684 0.970197
R1706 VGND.n714 VGND.n713 0.970197
R1707 VGND.n704 VGND.n683 0.970197
R1708 VGND.n803 VGND.n790 0.970197
R1709 VGND.n804 VGND.n789 0.970197
R1710 VGND.n798 VGND.n797 0.970197
R1711 VGND.n991 VGND.n954 0.970197
R1712 VGND.n998 VGND.n997 0.970197
R1713 VGND.n988 VGND.n953 0.970197
R1714 VGND.n928 VGND.n891 0.970197
R1715 VGND.n935 VGND.n934 0.970197
R1716 VGND.n925 VGND.n890 0.970197
R1717 VGND.n314 VGND.n301 0.970197
R1718 VGND.n315 VGND.n300 0.970197
R1719 VGND.n309 VGND.n308 0.970197
R1720 VGND.n423 VGND.n386 0.970197
R1721 VGND.n430 VGND.n429 0.970197
R1722 VGND.n420 VGND.n385 0.970197
R1723 VGND.n223 VGND.n221 0.927299
R1724 VGND.n471 VGND.n469 0.927299
R1725 VGND.n700 VGND.n698 0.927299
R1726 VGND.n786 VGND.n784 0.927299
R1727 VGND.n984 VGND.n982 0.927299
R1728 VGND.n921 VGND.n919 0.927299
R1729 VGND.n297 VGND.n295 0.927299
R1730 VGND.n416 VGND.n414 0.927299
R1731 VGND.n1066 VGND.n1 0.8465
R1732 VGND.n1067 VGND.n1066 0.8465
R1733 VGND.n249 VGND.n248 0.846456
R1734 VGND.n436 VGND.n78 0.846456
R1735 VGND.n820 VGND.n819 0.846456
R1736 VGND.n949 VGND.n948 0.846456
R1737 VGND.n1050 VGND.n1049 0.846456
R1738 VGND.n323 VGND.n322 0.846456
R1739 VGND.n381 VGND.n380 0.846456
R1740 VGND.n613 VGND.n566 0.721167
R1741 VGND.n209 VGND.n207 0.690273
R1742 VGND.n456 VGND.n454 0.690273
R1743 VGND.n679 VGND.n677 0.690273
R1744 VGND.n772 VGND.n770 0.690273
R1745 VGND.n969 VGND.n967 0.690273
R1746 VGND.n906 VGND.n904 0.690273
R1747 VGND.n283 VGND.n281 0.690273
R1748 VGND.n401 VGND.n399 0.690273
R1749 VGND.n221 VGND.n210 0.60675
R1750 VGND.n469 VGND.n458 0.60675
R1751 VGND.n698 VGND.n687 0.60675
R1752 VGND.n784 VGND.n773 0.60675
R1753 VGND.n982 VGND.n971 0.60675
R1754 VGND.n919 VGND.n908 0.60675
R1755 VGND.n295 VGND.n284 0.60675
R1756 VGND.n414 VGND.n403 0.60675
R1757 VGND.n1037 VGND.n59 0.5455
R1758 VGND.n719 VGND.n612 0.5455
R1759 VGND.n1004 VGND.n1003 0.5455
R1760 VGND.n940 VGND.n834 0.5455
R1761 VGND.n757 VGND.n756 0.5455
R1762 VGND.n518 VGND.n517 0.5455
R1763 VGND.n354 VGND.n0 0.5455
R1764 VGND.n1065 VGND.n1064 0.5455
R1765 VGND.n221 VGND.n215 0.516045
R1766 VGND.n469 VGND.n463 0.516045
R1767 VGND.n698 VGND.n692 0.516045
R1768 VGND.n784 VGND.n778 0.516045
R1769 VGND.n982 VGND.n976 0.516045
R1770 VGND.n919 VGND.n913 0.516045
R1771 VGND.n295 VGND.n289 0.516045
R1772 VGND.n414 VGND.n408 0.516045
R1773 VGND.n211 VGND.n210 0.454213
R1774 VGND.n459 VGND.n458 0.454213
R1775 VGND.n688 VGND.n687 0.454213
R1776 VGND.n774 VGND.n773 0.454213
R1777 VGND.n972 VGND.n971 0.454213
R1778 VGND.n909 VGND.n908 0.454213
R1779 VGND.n285 VGND.n284 0.454213
R1780 VGND.n404 VGND.n403 0.454213
R1781 VGND.n238 VGND.n237 0.363
R1782 VGND.n487 VGND.n486 0.363
R1783 VGND.n716 VGND.n715 0.363
R1784 VGND.n801 VGND.n800 0.363
R1785 VGND.n1000 VGND.n999 0.363
R1786 VGND.n937 VGND.n936 0.363
R1787 VGND.n312 VGND.n311 0.363
R1788 VGND.n432 VGND.n431 0.363
R1789 VGND.n218 VGND.n210 0.347226
R1790 VGND.n466 VGND.n458 0.347226
R1791 VGND.n695 VGND.n687 0.347226
R1792 VGND.n781 VGND.n773 0.347226
R1793 VGND.n979 VGND.n971 0.347226
R1794 VGND.n916 VGND.n908 0.347226
R1795 VGND.n292 VGND.n284 0.347226
R1796 VGND.n411 VGND.n403 0.347226
R1797 VGND.n236 VGND.n235 0.344944
R1798 VGND.n240 VGND.n239 0.344944
R1799 VGND.n440 VGND.n438 0.344944
R1800 VGND.n441 VGND.n439 0.344944
R1801 VGND.n683 VGND.n681 0.344944
R1802 VGND.n684 VGND.n682 0.344944
R1803 VGND.n799 VGND.n798 0.344944
R1804 VGND.n803 VGND.n802 0.344944
R1805 VGND.n953 VGND.n951 0.344944
R1806 VGND.n954 VGND.n952 0.344944
R1807 VGND.n890 VGND.n888 0.344944
R1808 VGND.n891 VGND.n889 0.344944
R1809 VGND.n310 VGND.n309 0.344944
R1810 VGND.n314 VGND.n313 0.344944
R1811 VGND.n385 VGND.n383 0.344944
R1812 VGND.n386 VGND.n384 0.344944
R1813 VGND.n212 VGND.n211 0.319807
R1814 VGND.n460 VGND.n459 0.319807
R1815 VGND.n689 VGND.n688 0.319807
R1816 VGND.n775 VGND.n774 0.319807
R1817 VGND.n973 VGND.n972 0.319807
R1818 VGND.n910 VGND.n909 0.319807
R1819 VGND.n286 VGND.n285 0.319807
R1820 VGND.n405 VGND.n404 0.319807
R1821 VGND.n215 VGND.n214 0.291342
R1822 VGND.n463 VGND.n462 0.291342
R1823 VGND.n692 VGND.n691 0.291342
R1824 VGND.n778 VGND.n777 0.291342
R1825 VGND.n976 VGND.n975 0.291342
R1826 VGND.n913 VGND.n912 0.291342
R1827 VGND.n289 VGND.n288 0.291342
R1828 VGND.n408 VGND.n407 0.291342
R1829 VGND.n218 VGND.n215 0.22669
R1830 VGND.n466 VGND.n463 0.22669
R1831 VGND.n695 VGND.n692 0.22669
R1832 VGND.n781 VGND.n778 0.22669
R1833 VGND.n979 VGND.n976 0.22669
R1834 VGND.n916 VGND.n913 0.22669
R1835 VGND.n292 VGND.n289 0.22669
R1836 VGND.n411 VGND.n408 0.22669
R1837 VGND.n246 VGND.n209 0.216409
R1838 VGND.n457 VGND.n456 0.216409
R1839 VGND.n680 VGND.n679 0.216409
R1840 VGND.n809 VGND.n772 0.216409
R1841 VGND.n970 VGND.n969 0.216409
R1842 VGND.n907 VGND.n906 0.216409
R1843 VGND.n320 VGND.n283 0.216409
R1844 VGND.n402 VGND.n401 0.216409
R1845 VGND.n245 VGND.n223 0.210727
R1846 VGND.n472 VGND.n471 0.210727
R1847 VGND.n701 VGND.n700 0.210727
R1848 VGND.n808 VGND.n786 0.210727
R1849 VGND.n985 VGND.n984 0.210727
R1850 VGND.n922 VGND.n921 0.210727
R1851 VGND.n319 VGND.n297 0.210727
R1852 VGND.n417 VGND.n416 0.210727
R1853 VGND VGND.n1069 0.198859
R1854 VGND.n248 VGND.n247 0.158833
R1855 VGND.n437 VGND.n436 0.158833
R1856 VGND.n820 VGND.n810 0.158833
R1857 VGND.n950 VGND.n949 0.158833
R1858 VGND.n1050 VGND.n41 0.158833
R1859 VGND.n322 VGND.n321 0.158833
R1860 VGND.n382 VGND.n381 0.158833
R1861 VGND.n216 VGND.n215 0.158238
R1862 VGND.n464 VGND.n463 0.158238
R1863 VGND.n693 VGND.n692 0.158238
R1864 VGND.n779 VGND.n778 0.158238
R1865 VGND.n977 VGND.n976 0.158238
R1866 VGND.n914 VGND.n913 0.158238
R1867 VGND.n290 VGND.n289 0.158238
R1868 VGND.n409 VGND.n408 0.158238
R1869 VGND.n517 VGND 0.149613
R1870 VGND VGND.n1065 0.14291
R1871 VGND.n516 VGND.n490 0.142507
R1872 VGND.n268 VGND.n27 0.142507
R1873 VGND.n194 VGND.n193 0.142507
R1874 VGND.n435 VGND.n121 0.1417
R1875 VGND.n233 VGND.n228 0.135283
R1876 VGND.n238 VGND.n226 0.135283
R1877 VGND.n477 VGND.n476 0.135283
R1878 VGND.n486 VGND.n485 0.135283
R1879 VGND.n706 VGND.n705 0.135283
R1880 VGND.n715 VGND.n714 0.135283
R1881 VGND.n796 VGND.n791 0.135283
R1882 VGND.n801 VGND.n789 0.135283
R1883 VGND.n990 VGND.n989 0.135283
R1884 VGND.n999 VGND.n998 0.135283
R1885 VGND.n927 VGND.n926 0.135283
R1886 VGND.n936 VGND.n935 0.135283
R1887 VGND.n307 VGND.n302 0.135283
R1888 VGND.n312 VGND.n300 0.135283
R1889 VGND.n422 VGND.n421 0.135283
R1890 VGND.n431 VGND.n430 0.135283
R1891 VGND VGND.n59 0.133711
R1892 VGND.n173 VGND.n172 0.120292
R1893 VGND.n173 VGND.n168 0.120292
R1894 VGND.n191 VGND.n169 0.120292
R1895 VGND.n186 VGND.n169 0.120292
R1896 VGND.n186 VGND.n185 0.120292
R1897 VGND.n185 VGND.n180 0.120292
R1898 VGND.n181 VGND.n180 0.120292
R1899 VGND.n101 VGND.n100 0.120292
R1900 VGND.n101 VGND.n96 0.120292
R1901 VGND.n119 VGND.n97 0.120292
R1902 VGND.n114 VGND.n97 0.120292
R1903 VGND.n114 VGND.n113 0.120292
R1904 VGND.n113 VGND.n108 0.120292
R1905 VGND.n109 VGND.n108 0.120292
R1906 VGND.n620 VGND.n619 0.120292
R1907 VGND.n620 VGND.n614 0.120292
R1908 VGND.n638 VGND.n615 0.120292
R1909 VGND.n633 VGND.n615 0.120292
R1910 VGND.n633 VGND.n632 0.120292
R1911 VGND.n632 VGND.n627 0.120292
R1912 VGND.n628 VGND.n627 0.120292
R1913 VGND.n646 VGND.n645 0.120292
R1914 VGND.n646 VGND.n641 0.120292
R1915 VGND.n664 VGND.n642 0.120292
R1916 VGND.n659 VGND.n642 0.120292
R1917 VGND.n659 VGND.n658 0.120292
R1918 VGND.n658 VGND.n653 0.120292
R1919 VGND.n654 VGND.n653 0.120292
R1920 VGND.n867 VGND.n866 0.120292
R1921 VGND.n867 VGND.n861 0.120292
R1922 VGND.n885 VGND.n862 0.120292
R1923 VGND.n880 VGND.n862 0.120292
R1924 VGND.n880 VGND.n879 0.120292
R1925 VGND.n879 VGND.n874 0.120292
R1926 VGND.n875 VGND.n874 0.120292
R1927 VGND.n840 VGND.n839 0.120292
R1928 VGND.n840 VGND.n835 0.120292
R1929 VGND.n858 VGND.n836 0.120292
R1930 VGND.n853 VGND.n836 0.120292
R1931 VGND.n853 VGND.n852 0.120292
R1932 VGND.n852 VGND.n847 0.120292
R1933 VGND.n848 VGND.n847 0.120292
R1934 VGND.n496 VGND.n495 0.120292
R1935 VGND.n496 VGND.n491 0.120292
R1936 VGND.n514 VGND.n492 0.120292
R1937 VGND.n509 VGND.n492 0.120292
R1938 VGND.n509 VGND.n508 0.120292
R1939 VGND.n508 VGND.n503 0.120292
R1940 VGND.n504 VGND.n503 0.120292
R1941 VGND.n7 VGND.n6 0.120292
R1942 VGND.n7 VGND.n2 0.120292
R1943 VGND.n25 VGND.n3 0.120292
R1944 VGND.n20 VGND.n3 0.120292
R1945 VGND.n20 VGND.n19 0.120292
R1946 VGND.n19 VGND.n14 0.120292
R1947 VGND.n15 VGND.n14 0.120292
R1948 VGND.n192 VGND.n168 0.112479
R1949 VGND.n120 VGND.n96 0.112479
R1950 VGND.n639 VGND.n614 0.112479
R1951 VGND.n665 VGND.n641 0.112479
R1952 VGND.n886 VGND.n861 0.112479
R1953 VGND.n859 VGND.n835 0.112479
R1954 VGND.n515 VGND.n491 0.112479
R1955 VGND.n26 VGND.n2 0.112479
R1956 VGND.n717 VGND.n680 0.0961731
R1957 VGND.n247 VGND.n246 0.09425
R1958 VGND.n457 VGND.n437 0.09425
R1959 VGND.n810 VGND.n809 0.09425
R1960 VGND.n970 VGND.n950 0.09425
R1961 VGND.n907 VGND.n41 0.09425
R1962 VGND.n321 VGND.n320 0.09425
R1963 VGND.n402 VGND.n382 0.09425
R1964 VGND.n490 VGND 0.0941643
R1965 VGND.n268 VGND 0.0941643
R1966 VGND.n194 VGND 0.0941643
R1967 VGND VGND.n435 0.0936321
R1968 VGND.n214 VGND.n213 0.0714406
R1969 VGND.n462 VGND.n461 0.0714406
R1970 VGND.n691 VGND.n690 0.0714406
R1971 VGND.n777 VGND.n776 0.0714406
R1972 VGND.n975 VGND.n974 0.0714406
R1973 VGND.n912 VGND.n911 0.0714406
R1974 VGND.n288 VGND.n287 0.0714406
R1975 VGND.n407 VGND.n406 0.0714406
R1976 VGND.n613 VGND 0.0610165
R1977 VGND.n172 VGND 0.0603958
R1978 VGND.n100 VGND 0.0603958
R1979 VGND.n619 VGND 0.0603958
R1980 VGND.n645 VGND 0.0603958
R1981 VGND.n866 VGND 0.0603958
R1982 VGND.n839 VGND 0.0603958
R1983 VGND.n495 VGND 0.0603958
R1984 VGND.n6 VGND 0.0603958
R1985 VGND.n717 VGND.n716 0.0599231
R1986 VGND.n196 VGND.n195 0.0584812
R1987 VGND.n489 VGND.n488 0.0584812
R1988 VGND.n718 VGND.n717 0.0584812
R1989 VGND.n759 VGND.n758 0.0584812
R1990 VGND.n1002 VGND.n1001 0.0584812
R1991 VGND.n939 VGND.n938 0.0584812
R1992 VGND.n270 VGND.n269 0.0584812
R1993 VGND.n434 VGND.n433 0.0584812
R1994 VGND.n517 VGND.n516 0.0582429
R1995 VGND.n1065 VGND.n27 0.0582429
R1996 VGND.n193 VGND.n59 0.0582429
R1997 VGND.n121 VGND.n0 0.0579148
R1998 VGND.n195 VGND 0.0520484
R1999 VGND.n489 VGND 0.0520484
R2000 VGND.n718 VGND 0.0520484
R2001 VGND.n758 VGND 0.0520484
R2002 VGND.n1002 VGND 0.0520484
R2003 VGND.n939 VGND 0.0520484
R2004 VGND.n269 VGND 0.0520484
R2005 VGND.n434 VGND 0.0520484
R2006 VGND.n1 VGND 0.0503372
R2007 VGND VGND.n355 0.0459545
R2008 VGND VGND.n1038 0.0459545
R2009 VGND.n1036 VGND 0.0459545
R2010 VGND.n755 VGND 0.0459545
R2011 VGND.n602 VGND 0.0459545
R2012 VGND.n611 VGND 0.0459545
R2013 VGND.n565 VGND 0.0459545
R2014 VGND VGND.n1005 0.0459545
R2015 VGND VGND.n567 0.0459545
R2016 VGND.n833 VGND 0.0459545
R2017 VGND VGND.n720 0.0459545
R2018 VGND VGND.n28 0.0459545
R2019 VGND VGND.n95 0.0459545
R2020 VGND VGND.n519 0.0459545
R2021 VGND.n353 VGND 0.0459545
R2022 VGND.n1063 VGND 0.0459545
R2023 VGND.n237 VGND.n196 0.0455
R2024 VGND.n488 VGND.n487 0.0455
R2025 VGND.n800 VGND.n759 0.0455
R2026 VGND.n1001 VGND.n1000 0.0455
R2027 VGND.n938 VGND.n937 0.0455
R2028 VGND.n311 VGND.n270 0.0455
R2029 VGND.n433 VGND.n432 0.0455
R2030 VGND.n202 VGND.n198 0.0429342
R2031 VGND.n203 VGND.n202 0.0429342
R2032 VGND.n204 VGND.n203 0.0429342
R2033 VGND.n204 VGND.n197 0.0429342
R2034 VGND.n449 VGND.n445 0.0429342
R2035 VGND.n450 VGND.n449 0.0429342
R2036 VGND.n451 VGND.n450 0.0429342
R2037 VGND.n451 VGND.n444 0.0429342
R2038 VGND.n672 VGND.n668 0.0429342
R2039 VGND.n673 VGND.n672 0.0429342
R2040 VGND.n674 VGND.n673 0.0429342
R2041 VGND.n674 VGND.n667 0.0429342
R2042 VGND.n765 VGND.n761 0.0429342
R2043 VGND.n766 VGND.n765 0.0429342
R2044 VGND.n767 VGND.n766 0.0429342
R2045 VGND.n767 VGND.n760 0.0429342
R2046 VGND.n962 VGND.n958 0.0429342
R2047 VGND.n963 VGND.n962 0.0429342
R2048 VGND.n964 VGND.n963 0.0429342
R2049 VGND.n964 VGND.n957 0.0429342
R2050 VGND.n899 VGND.n895 0.0429342
R2051 VGND.n900 VGND.n899 0.0429342
R2052 VGND.n901 VGND.n900 0.0429342
R2053 VGND.n901 VGND.n894 0.0429342
R2054 VGND.n276 VGND.n272 0.0429342
R2055 VGND.n277 VGND.n276 0.0429342
R2056 VGND.n278 VGND.n277 0.0429342
R2057 VGND.n278 VGND.n271 0.0429342
R2058 VGND.n394 VGND.n390 0.0429342
R2059 VGND.n395 VGND.n394 0.0429342
R2060 VGND.n396 VGND.n395 0.0429342
R2061 VGND.n396 VGND.n389 0.0429342
R2062 VGND.n200 VGND.n199 0.0389615
R2063 VGND.n447 VGND.n446 0.0389615
R2064 VGND.n670 VGND.n669 0.0389615
R2065 VGND.n763 VGND.n762 0.0389615
R2066 VGND.n960 VGND.n959 0.0389615
R2067 VGND.n897 VGND.n896 0.0389615
R2068 VGND.n274 VGND.n273 0.0389615
R2069 VGND.n392 VGND.n391 0.0389615
R2070 VGND.n207 VGND.n197 0.0340526
R2071 VGND.n454 VGND.n444 0.0340526
R2072 VGND.n677 VGND.n667 0.0340526
R2073 VGND.n770 VGND.n760 0.0340526
R2074 VGND.n967 VGND.n957 0.0340526
R2075 VGND.n904 VGND.n894 0.0340526
R2076 VGND.n281 VGND.n271 0.0340526
R2077 VGND.n399 VGND.n389 0.0340526
R2078 VGND.n355 VGND 0.0338333
R2079 VGND.n1038 VGND 0.0338333
R2080 VGND.n1036 VGND 0.0338333
R2081 VGND.n755 VGND 0.0338333
R2082 VGND.n602 VGND 0.0338333
R2083 VGND.n611 VGND 0.0338333
R2084 VGND.n565 VGND 0.0338333
R2085 VGND.n1005 VGND 0.0338333
R2086 VGND.n567 VGND 0.0338333
R2087 VGND.n833 VGND 0.0338333
R2088 VGND.n720 VGND 0.0338333
R2089 VGND.n28 VGND 0.0338333
R2090 VGND.n95 VGND 0.0338333
R2091 VGND.n519 VGND 0.0338333
R2092 VGND.n353 VGND 0.0338333
R2093 VGND.n1063 VGND 0.0338333
R2094 VGND.n215 VGND.n212 0.0289653
R2095 VGND.n463 VGND.n460 0.0289653
R2096 VGND.n692 VGND.n689 0.0289653
R2097 VGND.n778 VGND.n775 0.0289653
R2098 VGND.n976 VGND.n973 0.0289653
R2099 VGND.n913 VGND.n910 0.0289653
R2100 VGND.n289 VGND.n286 0.0289653
R2101 VGND.n408 VGND.n405 0.0289653
R2102 VGND.n1068 VGND.n0 0.0265369
R2103 VGND.n181 VGND 0.0226354
R2104 VGND.n109 VGND 0.0226354
R2105 VGND.n628 VGND 0.0226354
R2106 VGND.n654 VGND 0.0226354
R2107 VGND.n875 VGND 0.0226354
R2108 VGND.n848 VGND 0.0226354
R2109 VGND.n504 VGND 0.0226354
R2110 VGND.n15 VGND 0.0226354
R2111 VGND.n1068 VGND.n1067 0.0101424
R2112 VGND.n1069 VGND.n1068 0.0101424
R2113 VGND.n192 VGND.n191 0.0083125
R2114 VGND.n120 VGND.n119 0.0083125
R2115 VGND.n639 VGND.n638 0.0083125
R2116 VGND.n665 VGND.n664 0.0083125
R2117 VGND.n886 VGND.n885 0.0083125
R2118 VGND.n859 VGND.n858 0.0083125
R2119 VGND.n515 VGND.n514 0.0083125
R2120 VGND.n26 VGND.n25 0.0083125
R2121 VGND.n200 VGND.n198 0.00773684
R2122 VGND.n447 VGND.n445 0.00773684
R2123 VGND.n670 VGND.n668 0.00773684
R2124 VGND.n763 VGND.n761 0.00773684
R2125 VGND.n960 VGND.n958 0.00773684
R2126 VGND.n897 VGND.n895 0.00773684
R2127 VGND.n274 VGND.n272 0.00773684
R2128 VGND.n392 VGND.n390 0.00773684
R2129 VGND.n246 VGND.n245 0.00618182
R2130 VGND.n472 VGND.n457 0.00618182
R2131 VGND.n701 VGND.n680 0.00618182
R2132 VGND.n809 VGND.n808 0.00618182
R2133 VGND.n985 VGND.n970 0.00618182
R2134 VGND.n922 VGND.n907 0.00618182
R2135 VGND.n320 VGND.n319 0.00618182
R2136 VGND.n417 VGND.n402 0.00618182
R2137 VGND.n1066 VGND 0.00553571
R2138 VGND.n940 VGND.n939 0.00544203
R2139 VGND.n1003 VGND.n1002 0.00544203
R2140 VGND.n758 VGND.n757 0.00544203
R2141 VGND.n719 VGND.n718 0.00544203
R2142 VGND.n490 VGND.n489 0.00544203
R2143 VGND.n435 VGND.n434 0.00544203
R2144 VGND.n269 VGND.n268 0.00544203
R2145 VGND.n195 VGND.n194 0.00544203
R2146 VGND.n1003 VGND.n566 0.00167117
R2147 VGND.n247 VGND.n196 0.00154167
R2148 VGND.n488 VGND.n437 0.00154167
R2149 VGND.n810 VGND.n759 0.00154167
R2150 VGND.n1001 VGND.n950 0.00154167
R2151 VGND.n938 VGND.n41 0.00154167
R2152 VGND.n321 VGND.n270 0.00154167
R2153 VGND.n433 VGND.n382 0.00154167
R2154 VGND VGND.n613 0.000959214
R2155 VGND VGND.n1 0.000955654
R2156 VGND.n940 VGND.n887 0.0008453
R2157 VGND.n719 VGND.n666 0.000770545
R2158 VGND.n757 VGND.n719 0.000710028
R2159 VGND.n666 VGND.n640 0.000710028
R2160 VGND.n1003 VGND.n940 0.000635272
R2161 VGND.n887 VGND.n860 0.000635272
R2162 VGND.n860 VGND 0.000613914
R2163 VGND.n640 VGND 0.000539158
R2164 VPWR.n174 VPWR.n173 18810
R2165 VPWR.n253 VPWR.n252 18810
R2166 VPWR.n93 VPWR.n92 18810
R2167 VPWR.n14 VPWR.n13 18810
R2168 VPWR.n455 VPWR.n454 18810
R2169 VPWR.n374 VPWR.n373 18810
R2170 VPWR.n617 VPWR.n616 18810
R2171 VPWR.n536 VPWR.n535 18810
R2172 VPWR.n175 VPWR.n174 18786.2
R2173 VPWR.n175 VPWR.n166 18786.2
R2174 VPWR.n254 VPWR.n253 18786.2
R2175 VPWR.n254 VPWR.n245 18786.2
R2176 VPWR.n94 VPWR.n93 18786.2
R2177 VPWR.n94 VPWR.n85 18786.2
R2178 VPWR.n15 VPWR.n14 18786.2
R2179 VPWR.n15 VPWR.n6 18786.2
R2180 VPWR.n456 VPWR.n455 18786.2
R2181 VPWR.n456 VPWR.n447 18786.2
R2182 VPWR.n375 VPWR.n374 18786.2
R2183 VPWR.n375 VPWR.n366 18786.2
R2184 VPWR.n618 VPWR.n617 18786.2
R2185 VPWR.n618 VPWR.n609 18786.2
R2186 VPWR.n537 VPWR.n536 18786.2
R2187 VPWR.n537 VPWR.n528 18786.2
R2188 VPWR.n173 VPWR.n166 18667.5
R2189 VPWR.n252 VPWR.n245 18667.5
R2190 VPWR.n92 VPWR.n85 18667.5
R2191 VPWR.n13 VPWR.n6 18667.5
R2192 VPWR.n454 VPWR.n447 18667.5
R2193 VPWR.n373 VPWR.n366 18667.5
R2194 VPWR.n616 VPWR.n609 18667.5
R2195 VPWR.n535 VPWR.n528 18667.5
R2196 VPWR.n176 VPWR.n164 7334.54
R2197 VPWR.n255 VPWR.n243 7334.54
R2198 VPWR.n95 VPWR.n83 7334.54
R2199 VPWR.n16 VPWR.n4 7334.54
R2200 VPWR.n457 VPWR.n445 7334.54
R2201 VPWR.n376 VPWR.n364 7334.54
R2202 VPWR.n619 VPWR.n607 7334.54
R2203 VPWR.n538 VPWR.n526 7334.54
R2204 VPWR.n172 VPWR.n165 7332.73
R2205 VPWR.n251 VPWR.n244 7332.73
R2206 VPWR.n91 VPWR.n84 7332.73
R2207 VPWR.n12 VPWR.n5 7332.73
R2208 VPWR.n453 VPWR.n446 7332.73
R2209 VPWR.n372 VPWR.n365 7332.73
R2210 VPWR.n615 VPWR.n608 7332.73
R2211 VPWR.n534 VPWR.n527 7332.73
R2212 VPWR.n176 VPWR.n165 7312.73
R2213 VPWR.n255 VPWR.n244 7312.73
R2214 VPWR.n95 VPWR.n84 7312.73
R2215 VPWR.n16 VPWR.n5 7312.73
R2216 VPWR.n457 VPWR.n446 7312.73
R2217 VPWR.n376 VPWR.n365 7312.73
R2218 VPWR.n619 VPWR.n608 7312.73
R2219 VPWR.n538 VPWR.n527 7312.73
R2220 VPWR.n172 VPWR.n164 7300
R2221 VPWR.n251 VPWR.n243 7300
R2222 VPWR.n91 VPWR.n83 7300
R2223 VPWR.n12 VPWR.n4 7300
R2224 VPWR.n453 VPWR.n445 7300
R2225 VPWR.n372 VPWR.n364 7300
R2226 VPWR.n615 VPWR.n607 7300
R2227 VPWR.n534 VPWR.n526 7300
R2228 VPWR.n227 VPWR.n225 4136.47
R2229 VPWR.n234 VPWR.n232 4136.47
R2230 VPWR.n306 VPWR.n304 4136.47
R2231 VPWR.n313 VPWR.n311 4136.47
R2232 VPWR.n67 VPWR.n65 4136.47
R2233 VPWR.n74 VPWR.n72 4136.47
R2234 VPWR.n146 VPWR.n144 4136.47
R2235 VPWR.n153 VPWR.n151 4136.47
R2236 VPWR.n403 VPWR.n401 4136.47
R2237 VPWR.n410 VPWR.n408 4136.47
R2238 VPWR.n323 VPWR.n321 4136.47
R2239 VPWR.n330 VPWR.n328 4136.47
R2240 VPWR.n565 VPWR.n563 4136.47
R2241 VPWR.n572 VPWR.n570 4136.47
R2242 VPWR.n485 VPWR.n483 4136.47
R2243 VPWR.n492 VPWR.n490 4136.47
R2244 VPWR.n227 VPWR.n224 2068.24
R2245 VPWR.n234 VPWR.n231 2068.24
R2246 VPWR.n306 VPWR.n303 2068.24
R2247 VPWR.n313 VPWR.n310 2068.24
R2248 VPWR.n67 VPWR.n64 2068.24
R2249 VPWR.n74 VPWR.n71 2068.24
R2250 VPWR.n146 VPWR.n143 2068.24
R2251 VPWR.n153 VPWR.n150 2068.24
R2252 VPWR.n403 VPWR.n400 2068.24
R2253 VPWR.n410 VPWR.n407 2068.24
R2254 VPWR.n323 VPWR.n320 2068.24
R2255 VPWR.n330 VPWR.n327 2068.24
R2256 VPWR.n565 VPWR.n562 2068.24
R2257 VPWR.n572 VPWR.n569 2068.24
R2258 VPWR.n485 VPWR.n482 2068.24
R2259 VPWR.n492 VPWR.n489 2068.24
R2260 VPWR.n170 VPWR.n168 781.188
R2261 VPWR.n249 VPWR.n247 781.188
R2262 VPWR.n89 VPWR.n87 781.188
R2263 VPWR.n10 VPWR.n8 781.188
R2264 VPWR.n451 VPWR.n449 781.188
R2265 VPWR.n370 VPWR.n368 781.188
R2266 VPWR.n613 VPWR.n611 781.188
R2267 VPWR.n532 VPWR.n530 781.188
R2268 VPWR.n178 VPWR.n162 779.442
R2269 VPWR.n257 VPWR.n241 779.442
R2270 VPWR.n97 VPWR.n81 779.442
R2271 VPWR.n18 VPWR.n2 779.442
R2272 VPWR.n459 VPWR.n443 779.442
R2273 VPWR.n378 VPWR.n362 779.442
R2274 VPWR.n621 VPWR.n605 779.442
R2275 VPWR.n540 VPWR.n524 779.442
R2276 VPWR.n177 VPWR.n163 779.056
R2277 VPWR.n256 VPWR.n242 779.056
R2278 VPWR.n96 VPWR.n82 779.056
R2279 VPWR.n17 VPWR.n3 779.056
R2280 VPWR.n458 VPWR.n444 779.056
R2281 VPWR.n377 VPWR.n363 779.056
R2282 VPWR.n620 VPWR.n606 779.056
R2283 VPWR.n539 VPWR.n525 779.056
R2284 VPWR.n171 VPWR.n167 778.668
R2285 VPWR.n250 VPWR.n246 778.668
R2286 VPWR.n90 VPWR.n86 778.668
R2287 VPWR.n11 VPWR.n7 778.668
R2288 VPWR.n452 VPWR.n448 778.668
R2289 VPWR.n371 VPWR.n367 778.668
R2290 VPWR.n614 VPWR.n610 778.668
R2291 VPWR.n533 VPWR.n529 778.668
R2292 VPWR.t298 VPWR.t254 478.712
R2293 VPWR.t304 VPWR.t298 478.712
R2294 VPWR.t308 VPWR.t304 478.712
R2295 VPWR.t296 VPWR.t308 478.712
R2296 VPWR.t294 VPWR.t296 478.712
R2297 VPWR.t300 VPWR.t302 478.712
R2298 VPWR.t302 VPWR.t306 478.712
R2299 VPWR.t306 VPWR.t292 478.712
R2300 VPWR.t292 VPWR.t310 478.712
R2301 VPWR.t310 VPWR.t248 478.712
R2302 VPWR.t141 VPWR.t236 478.712
R2303 VPWR.t145 VPWR.t141 478.712
R2304 VPWR.t151 VPWR.t145 478.712
R2305 VPWR.t137 VPWR.t151 478.712
R2306 VPWR.t155 VPWR.t137 478.712
R2307 VPWR.t139 VPWR.t143 478.712
R2308 VPWR.t143 VPWR.t149 478.712
R2309 VPWR.t149 VPWR.t147 478.712
R2310 VPWR.t147 VPWR.t153 478.712
R2311 VPWR.t153 VPWR.t242 478.712
R2312 VPWR.t212 VPWR.t251 478.712
R2313 VPWR.t222 VPWR.t212 478.712
R2314 VPWR.t226 VPWR.t222 478.712
R2315 VPWR.t210 VPWR.t226 478.712
R2316 VPWR.t218 VPWR.t210 478.712
R2317 VPWR.t216 VPWR.t220 478.712
R2318 VPWR.t220 VPWR.t224 478.712
R2319 VPWR.t224 VPWR.t208 478.712
R2320 VPWR.t208 VPWR.t214 478.712
R2321 VPWR.t214 VPWR.t245 478.712
R2322 VPWR.t73 VPWR.t266 478.712
R2323 VPWR.t57 VPWR.t73 478.712
R2324 VPWR.t61 VPWR.t57 478.712
R2325 VPWR.t65 VPWR.t61 478.712
R2326 VPWR.t69 VPWR.t65 478.712
R2327 VPWR.t71 VPWR.t75 478.712
R2328 VPWR.t75 VPWR.t59 478.712
R2329 VPWR.t59 VPWR.t63 478.712
R2330 VPWR.t63 VPWR.t67 478.712
R2331 VPWR.t67 VPWR.t260 478.712
R2332 VPWR.t23 VPWR.t230 478.712
R2333 VPWR.t27 VPWR.t23 478.712
R2334 VPWR.t31 VPWR.t27 478.712
R2335 VPWR.t19 VPWR.t31 478.712
R2336 VPWR.t17 VPWR.t19 478.712
R2337 VPWR.t25 VPWR.t21 478.712
R2338 VPWR.t21 VPWR.t29 478.712
R2339 VPWR.t29 VPWR.t15 478.712
R2340 VPWR.t15 VPWR.t13 478.712
R2341 VPWR.t13 VPWR.t257 478.712
R2342 VPWR.t194 VPWR.t233 478.712
R2343 VPWR.t192 VPWR.t194 478.712
R2344 VPWR.t198 VPWR.t192 478.712
R2345 VPWR.t186 VPWR.t198 478.712
R2346 VPWR.t204 VPWR.t186 478.712
R2347 VPWR.t190 VPWR.t188 478.712
R2348 VPWR.t188 VPWR.t196 478.712
R2349 VPWR.t196 VPWR.t200 478.712
R2350 VPWR.t200 VPWR.t202 478.712
R2351 VPWR.t202 VPWR.t239 478.712
R2352 VPWR.t129 VPWR.t275 478.712
R2353 VPWR.t119 VPWR.t129 478.712
R2354 VPWR.t117 VPWR.t119 478.712
R2355 VPWR.t123 VPWR.t117 478.712
R2356 VPWR.t127 VPWR.t123 478.712
R2357 VPWR.t131 VPWR.t115 478.712
R2358 VPWR.t115 VPWR.t113 478.712
R2359 VPWR.t113 VPWR.t121 478.712
R2360 VPWR.t121 VPWR.t125 478.712
R2361 VPWR.t125 VPWR.t272 478.712
R2362 VPWR.t181 VPWR.t269 478.712
R2363 VPWR.t167 VPWR.t181 478.712
R2364 VPWR.t169 VPWR.t167 478.712
R2365 VPWR.t173 VPWR.t169 478.712
R2366 VPWR.t179 VPWR.t173 478.712
R2367 VPWR.t177 VPWR.t165 478.712
R2368 VPWR.t165 VPWR.t183 478.712
R2369 VPWR.t183 VPWR.t171 478.712
R2370 VPWR.t171 VPWR.t175 478.712
R2371 VPWR.t175 VPWR.t263 478.712
R2372 VPWR.n227 VPWR.t54 452.676
R2373 VPWR.t35 VPWR.n225 452.676
R2374 VPWR.n234 VPWR.t280 452.676
R2375 VPWR.t279 VPWR.n232 452.676
R2376 VPWR.n306 VPWR.t278 452.676
R2377 VPWR.t158 VPWR.n304 452.676
R2378 VPWR.n313 VPWR.t207 452.676
R2379 VPWR.t206 VPWR.n311 452.676
R2380 VPWR.n67 VPWR.t287 452.676
R2381 VPWR.t46 VPWR.n65 452.676
R2382 VPWR.n74 VPWR.t98 452.676
R2383 VPWR.t97 VPWR.n72 452.676
R2384 VPWR.n146 VPWR.t88 452.676
R2385 VPWR.t105 VPWR.n144 452.676
R2386 VPWR.n153 VPWR.t79 452.676
R2387 VPWR.t78 VPWR.n151 452.676
R2388 VPWR.n403 VPWR.t0 452.676
R2389 VPWR.t8 VPWR.n401 452.676
R2390 VPWR.n410 VPWR.t52 452.676
R2391 VPWR.t53 VPWR.n408 452.676
R2392 VPWR.n323 VPWR.t134 452.676
R2393 VPWR.t289 VPWR.n321 452.676
R2394 VPWR.n330 VPWR.t56 452.676
R2395 VPWR.t55 VPWR.n328 452.676
R2396 VPWR.n565 VPWR.t40 452.676
R2397 VPWR.t284 VPWR.n563 452.676
R2398 VPWR.n572 VPWR.t164 452.676
R2399 VPWR.t163 VPWR.n570 452.676
R2400 VPWR.n485 VPWR.t77 452.676
R2401 VPWR.t90 VPWR.n483 452.676
R2402 VPWR.n492 VPWR.t286 452.676
R2403 VPWR.t285 VPWR.n490 452.676
R2404 VPWR.n213 VPWR.t101 342.377
R2405 VPWR.n292 VPWR.t161 342.377
R2406 VPWR.n132 VPWR.t86 342.377
R2407 VPWR.n53 VPWR.t48 342.377
R2408 VPWR.n430 VPWR.t2 342.377
R2409 VPWR.n349 VPWR.t291 342.377
R2410 VPWR.n592 VPWR.t39 342.377
R2411 VPWR.n511 VPWR.t91 342.377
R2412 VPWR.n203 VPWR.t81 338.892
R2413 VPWR.n282 VPWR.t38 338.892
R2414 VPWR.n122 VPWR.t104 338.892
R2415 VPWR.n43 VPWR.t111 338.892
R2416 VPWR.n420 VPWR.t5 338.892
R2417 VPWR.n339 VPWR.t136 338.892
R2418 VPWR.n582 VPWR.t282 338.892
R2419 VPWR.n501 VPWR.t82 338.892
R2420 VPWR.n218 VPWR.n211 320.976
R2421 VPWR.n210 VPWR.n200 320.976
R2422 VPWR.n208 VPWR.n201 320.976
R2423 VPWR.n297 VPWR.n290 320.976
R2424 VPWR.n289 VPWR.n279 320.976
R2425 VPWR.n287 VPWR.n280 320.976
R2426 VPWR.n137 VPWR.n130 320.976
R2427 VPWR.n129 VPWR.n119 320.976
R2428 VPWR.n127 VPWR.n120 320.976
R2429 VPWR.n58 VPWR.n51 320.976
R2430 VPWR.n50 VPWR.n40 320.976
R2431 VPWR.n48 VPWR.n41 320.976
R2432 VPWR.n435 VPWR.n428 320.976
R2433 VPWR.n427 VPWR.n417 320.976
R2434 VPWR.n425 VPWR.n418 320.976
R2435 VPWR.n354 VPWR.n347 320.976
R2436 VPWR.n346 VPWR.n336 320.976
R2437 VPWR.n344 VPWR.n337 320.976
R2438 VPWR.n597 VPWR.n590 320.976
R2439 VPWR.n589 VPWR.n579 320.976
R2440 VPWR.n587 VPWR.n580 320.976
R2441 VPWR.n516 VPWR.n509 320.976
R2442 VPWR.n508 VPWR.n498 320.976
R2443 VPWR.n506 VPWR.n499 320.976
R2444 VPWR.n192 VPWR.t95 269.151
R2445 VPWR.n271 VPWR.t108 269.151
R2446 VPWR.n111 VPWR.t106 269.151
R2447 VPWR.n32 VPWR.t107 269.151
R2448 VPWR.n473 VPWR.t51 269.151
R2449 VPWR.n392 VPWR.t277 269.151
R2450 VPWR.n635 VPWR.t41 269.151
R2451 VPWR.n554 VPWR.t162 269.151
R2452 VPWR.n191 VPWR.t300 269.043
R2453 VPWR.n270 VPWR.t139 269.043
R2454 VPWR.n110 VPWR.t216 269.043
R2455 VPWR.n31 VPWR.t71 269.043
R2456 VPWR.n472 VPWR.t25 269.043
R2457 VPWR.n391 VPWR.t190 269.043
R2458 VPWR.n634 VPWR.t131 269.043
R2459 VPWR.n553 VPWR.t177 269.043
R2460 VPWR.n186 VPWR.t249 228.215
R2461 VPWR.n181 VPWR.t255 228.215
R2462 VPWR.n265 VPWR.t243 228.215
R2463 VPWR.n260 VPWR.t237 228.215
R2464 VPWR.n105 VPWR.t246 228.215
R2465 VPWR.n100 VPWR.t252 228.215
R2466 VPWR.n26 VPWR.t261 228.215
R2467 VPWR.n21 VPWR.t267 228.215
R2468 VPWR.n467 VPWR.t258 228.215
R2469 VPWR.n462 VPWR.t231 228.215
R2470 VPWR.n386 VPWR.t240 228.215
R2471 VPWR.n381 VPWR.t234 228.215
R2472 VPWR.n629 VPWR.t273 228.215
R2473 VPWR.n624 VPWR.t276 228.215
R2474 VPWR.n548 VPWR.t264 228.215
R2475 VPWR.n543 VPWR.t270 228.215
R2476 VPWR.t54 VPWR.n226 215.757
R2477 VPWR.n226 VPWR.t35 215.757
R2478 VPWR.t280 VPWR.n233 215.757
R2479 VPWR.n233 VPWR.t279 215.757
R2480 VPWR.t278 VPWR.n305 215.757
R2481 VPWR.n305 VPWR.t158 215.757
R2482 VPWR.t207 VPWR.n312 215.757
R2483 VPWR.n312 VPWR.t206 215.757
R2484 VPWR.t287 VPWR.n66 215.757
R2485 VPWR.n66 VPWR.t46 215.757
R2486 VPWR.t98 VPWR.n73 215.757
R2487 VPWR.n73 VPWR.t97 215.757
R2488 VPWR.t88 VPWR.n145 215.757
R2489 VPWR.n145 VPWR.t105 215.757
R2490 VPWR.t79 VPWR.n152 215.757
R2491 VPWR.n152 VPWR.t78 215.757
R2492 VPWR.t0 VPWR.n402 215.757
R2493 VPWR.n402 VPWR.t8 215.757
R2494 VPWR.t52 VPWR.n409 215.757
R2495 VPWR.n409 VPWR.t53 215.757
R2496 VPWR.t134 VPWR.n322 215.757
R2497 VPWR.n322 VPWR.t289 215.757
R2498 VPWR.t56 VPWR.n329 215.757
R2499 VPWR.n329 VPWR.t55 215.757
R2500 VPWR.t40 VPWR.n564 215.757
R2501 VPWR.n564 VPWR.t284 215.757
R2502 VPWR.t164 VPWR.n571 215.757
R2503 VPWR.n571 VPWR.t163 215.757
R2504 VPWR.t77 VPWR.n484 215.757
R2505 VPWR.n484 VPWR.t90 215.757
R2506 VPWR.t286 VPWR.n491 215.757
R2507 VPWR.n491 VPWR.t285 215.757
R2508 VPWR.n191 VPWR.t294 209.668
R2509 VPWR.n270 VPWR.t155 209.668
R2510 VPWR.n110 VPWR.t218 209.668
R2511 VPWR.n31 VPWR.t69 209.668
R2512 VPWR.n472 VPWR.t17 209.668
R2513 VPWR.n391 VPWR.t204 209.668
R2514 VPWR.n634 VPWR.t127 209.668
R2515 VPWR.n553 VPWR.t179 209.668
R2516 VPWR.n188 VPWR.n187 199.851
R2517 VPWR.n190 VPWR.n189 199.851
R2518 VPWR.n183 VPWR.n182 199.851
R2519 VPWR.n185 VPWR.n184 199.851
R2520 VPWR.n195 VPWR.n194 199.851
R2521 VPWR.n267 VPWR.n266 199.851
R2522 VPWR.n269 VPWR.n268 199.851
R2523 VPWR.n262 VPWR.n261 199.851
R2524 VPWR.n264 VPWR.n263 199.851
R2525 VPWR.n274 VPWR.n273 199.851
R2526 VPWR.n107 VPWR.n106 199.851
R2527 VPWR.n109 VPWR.n108 199.851
R2528 VPWR.n102 VPWR.n101 199.851
R2529 VPWR.n104 VPWR.n103 199.851
R2530 VPWR.n114 VPWR.n113 199.851
R2531 VPWR.n28 VPWR.n27 199.851
R2532 VPWR.n30 VPWR.n29 199.851
R2533 VPWR.n23 VPWR.n22 199.851
R2534 VPWR.n25 VPWR.n24 199.851
R2535 VPWR.n35 VPWR.n34 199.851
R2536 VPWR.n469 VPWR.n468 199.851
R2537 VPWR.n471 VPWR.n470 199.851
R2538 VPWR.n464 VPWR.n463 199.851
R2539 VPWR.n466 VPWR.n465 199.851
R2540 VPWR.n476 VPWR.n475 199.851
R2541 VPWR.n388 VPWR.n387 199.851
R2542 VPWR.n390 VPWR.n389 199.851
R2543 VPWR.n383 VPWR.n382 199.851
R2544 VPWR.n385 VPWR.n384 199.851
R2545 VPWR.n395 VPWR.n394 199.851
R2546 VPWR.n631 VPWR.n630 199.851
R2547 VPWR.n633 VPWR.n632 199.851
R2548 VPWR.n626 VPWR.n625 199.851
R2549 VPWR.n628 VPWR.n627 199.851
R2550 VPWR.n638 VPWR.n637 199.851
R2551 VPWR.n550 VPWR.n549 199.851
R2552 VPWR.n552 VPWR.n551 199.851
R2553 VPWR.n545 VPWR.n544 199.851
R2554 VPWR.n547 VPWR.n546 199.851
R2555 VPWR.n557 VPWR.n556 199.851
R2556 VPWR.n225 VPWR.n223 163.684
R2557 VPWR.n232 VPWR.n230 163.684
R2558 VPWR.n304 VPWR.n302 163.684
R2559 VPWR.n311 VPWR.n309 163.684
R2560 VPWR.n65 VPWR.n63 163.684
R2561 VPWR.n72 VPWR.n70 163.684
R2562 VPWR.n144 VPWR.n142 163.684
R2563 VPWR.n151 VPWR.n149 163.684
R2564 VPWR.n401 VPWR.n399 163.684
R2565 VPWR.n408 VPWR.n406 163.684
R2566 VPWR.n321 VPWR.n319 163.684
R2567 VPWR.n328 VPWR.n326 163.684
R2568 VPWR.n563 VPWR.n561 163.684
R2569 VPWR.n570 VPWR.n568 163.684
R2570 VPWR.n483 VPWR.n481 163.684
R2571 VPWR.n490 VPWR.n488 163.684
R2572 VPWR.n181 VPWR.t253 120.855
R2573 VPWR.n260 VPWR.t235 120.855
R2574 VPWR.n100 VPWR.t250 120.855
R2575 VPWR.n21 VPWR.t265 120.855
R2576 VPWR.n462 VPWR.t229 120.855
R2577 VPWR.n381 VPWR.t232 120.855
R2578 VPWR.n624 VPWR.t274 120.855
R2579 VPWR.n543 VPWR.t268 120.855
R2580 VPWR.n186 VPWR.t247 120.749
R2581 VPWR.n265 VPWR.t241 120.749
R2582 VPWR.n105 VPWR.t244 120.749
R2583 VPWR.n26 VPWR.t259 120.749
R2584 VPWR.n467 VPWR.t256 120.749
R2585 VPWR.n386 VPWR.t238 120.749
R2586 VPWR.n629 VPWR.t271 120.749
R2587 VPWR.n548 VPWR.t262 120.749
R2588 VPWR.n228 VPWR.n223 113.915
R2589 VPWR.n235 VPWR.n230 113.915
R2590 VPWR.n307 VPWR.n302 113.915
R2591 VPWR.n314 VPWR.n309 113.915
R2592 VPWR.n68 VPWR.n63 113.915
R2593 VPWR.n75 VPWR.n70 113.915
R2594 VPWR.n147 VPWR.n142 113.915
R2595 VPWR.n154 VPWR.n149 113.915
R2596 VPWR.n404 VPWR.n399 113.915
R2597 VPWR.n411 VPWR.n406 113.915
R2598 VPWR.n324 VPWR.n319 113.915
R2599 VPWR.n331 VPWR.n326 113.915
R2600 VPWR.n566 VPWR.n561 113.915
R2601 VPWR.n573 VPWR.n568 113.915
R2602 VPWR.n486 VPWR.n481 113.915
R2603 VPWR.n493 VPWR.n488 113.915
R2604 VPWR.n228 VPWR.n227 47.0382
R2605 VPWR.n235 VPWR.n234 47.0382
R2606 VPWR.n307 VPWR.n306 47.0382
R2607 VPWR.n314 VPWR.n313 47.0382
R2608 VPWR.n68 VPWR.n67 47.0382
R2609 VPWR.n75 VPWR.n74 47.0382
R2610 VPWR.n147 VPWR.n146 47.0382
R2611 VPWR.n154 VPWR.n153 47.0382
R2612 VPWR.n404 VPWR.n403 47.0382
R2613 VPWR.n411 VPWR.n410 47.0382
R2614 VPWR.n324 VPWR.n323 47.0382
R2615 VPWR.n331 VPWR.n330 47.0382
R2616 VPWR.n566 VPWR.n565 47.0382
R2617 VPWR.n573 VPWR.n572 47.0382
R2618 VPWR.n486 VPWR.n485 47.0382
R2619 VPWR.n493 VPWR.n492 47.0382
R2620 VPWR.n192 VPWR.n191 38.8096
R2621 VPWR.n271 VPWR.n270 38.8096
R2622 VPWR.n111 VPWR.n110 38.8096
R2623 VPWR.n32 VPWR.n31 38.8096
R2624 VPWR.n473 VPWR.n472 38.8096
R2625 VPWR.n392 VPWR.n391 38.8096
R2626 VPWR.n635 VPWR.n634 38.8096
R2627 VPWR.n554 VPWR.n553 38.8096
R2628 VPWR.n203 VPWR 35.5709
R2629 VPWR.n282 VPWR 35.5709
R2630 VPWR.n122 VPWR 35.5709
R2631 VPWR.n43 VPWR 35.5709
R2632 VPWR.n420 VPWR 35.5709
R2633 VPWR.n339 VPWR 35.5709
R2634 VPWR.n582 VPWR 35.5709
R2635 VPWR.n501 VPWR 35.5709
R2636 VPWR.n207 VPWR.n202 34.6358
R2637 VPWR.n220 VPWR.n219 34.6358
R2638 VPWR.n217 VPWR.n212 34.6358
R2639 VPWR.n286 VPWR.n281 34.6358
R2640 VPWR.n299 VPWR.n298 34.6358
R2641 VPWR.n296 VPWR.n291 34.6358
R2642 VPWR.n126 VPWR.n121 34.6358
R2643 VPWR.n139 VPWR.n138 34.6358
R2644 VPWR.n136 VPWR.n131 34.6358
R2645 VPWR.n47 VPWR.n42 34.6358
R2646 VPWR.n60 VPWR.n59 34.6358
R2647 VPWR.n57 VPWR.n52 34.6358
R2648 VPWR.n424 VPWR.n419 34.6358
R2649 VPWR.n437 VPWR.n436 34.6358
R2650 VPWR.n434 VPWR.n429 34.6358
R2651 VPWR.n343 VPWR.n338 34.6358
R2652 VPWR.n356 VPWR.n355 34.6358
R2653 VPWR.n353 VPWR.n348 34.6358
R2654 VPWR.n586 VPWR.n581 34.6358
R2655 VPWR.n599 VPWR.n598 34.6358
R2656 VPWR.n596 VPWR.n591 34.6358
R2657 VPWR.n505 VPWR.n500 34.6358
R2658 VPWR.n518 VPWR.n517 34.6358
R2659 VPWR.n515 VPWR.n510 34.6358
R2660 VPWR.n210 VPWR.n209 32.0005
R2661 VPWR.n289 VPWR.n288 32.0005
R2662 VPWR.n129 VPWR.n128 32.0005
R2663 VPWR.n50 VPWR.n49 32.0005
R2664 VPWR.n427 VPWR.n426 32.0005
R2665 VPWR.n346 VPWR.n345 32.0005
R2666 VPWR.n589 VPWR.n588 32.0005
R2667 VPWR.n508 VPWR.n507 32.0005
R2668 VPWR.n209 VPWR.n208 31.2476
R2669 VPWR.n288 VPWR.n287 31.2476
R2670 VPWR.n128 VPWR.n127 31.2476
R2671 VPWR.n49 VPWR.n48 31.2476
R2672 VPWR.n426 VPWR.n425 31.2476
R2673 VPWR.n345 VPWR.n344 31.2476
R2674 VPWR.n588 VPWR.n587 31.2476
R2675 VPWR.n507 VPWR.n506 31.2476
R2676 VPWR.n187 VPWR.t293 28.5655
R2677 VPWR.n187 VPWR.t311 28.5655
R2678 VPWR.n189 VPWR.t303 28.5655
R2679 VPWR.n189 VPWR.t307 28.5655
R2680 VPWR.n182 VPWR.t299 28.5655
R2681 VPWR.n182 VPWR.t305 28.5655
R2682 VPWR.n184 VPWR.t309 28.5655
R2683 VPWR.n184 VPWR.t297 28.5655
R2684 VPWR.n194 VPWR.t295 28.5655
R2685 VPWR.n194 VPWR.t301 28.5655
R2686 VPWR.n266 VPWR.t148 28.5655
R2687 VPWR.n266 VPWR.t154 28.5655
R2688 VPWR.n268 VPWR.t144 28.5655
R2689 VPWR.n268 VPWR.t150 28.5655
R2690 VPWR.n261 VPWR.t142 28.5655
R2691 VPWR.n261 VPWR.t146 28.5655
R2692 VPWR.n263 VPWR.t152 28.5655
R2693 VPWR.n263 VPWR.t138 28.5655
R2694 VPWR.n273 VPWR.t156 28.5655
R2695 VPWR.n273 VPWR.t140 28.5655
R2696 VPWR.n106 VPWR.t209 28.5655
R2697 VPWR.n106 VPWR.t215 28.5655
R2698 VPWR.n108 VPWR.t221 28.5655
R2699 VPWR.n108 VPWR.t225 28.5655
R2700 VPWR.n101 VPWR.t213 28.5655
R2701 VPWR.n101 VPWR.t223 28.5655
R2702 VPWR.n103 VPWR.t227 28.5655
R2703 VPWR.n103 VPWR.t211 28.5655
R2704 VPWR.n113 VPWR.t219 28.5655
R2705 VPWR.n113 VPWR.t217 28.5655
R2706 VPWR.n27 VPWR.t64 28.5655
R2707 VPWR.n27 VPWR.t68 28.5655
R2708 VPWR.n29 VPWR.t76 28.5655
R2709 VPWR.n29 VPWR.t60 28.5655
R2710 VPWR.n22 VPWR.t74 28.5655
R2711 VPWR.n22 VPWR.t58 28.5655
R2712 VPWR.n24 VPWR.t62 28.5655
R2713 VPWR.n24 VPWR.t66 28.5655
R2714 VPWR.n34 VPWR.t70 28.5655
R2715 VPWR.n34 VPWR.t72 28.5655
R2716 VPWR.n468 VPWR.t16 28.5655
R2717 VPWR.n468 VPWR.t14 28.5655
R2718 VPWR.n470 VPWR.t22 28.5655
R2719 VPWR.n470 VPWR.t30 28.5655
R2720 VPWR.n463 VPWR.t24 28.5655
R2721 VPWR.n463 VPWR.t28 28.5655
R2722 VPWR.n465 VPWR.t32 28.5655
R2723 VPWR.n465 VPWR.t20 28.5655
R2724 VPWR.n475 VPWR.t18 28.5655
R2725 VPWR.n475 VPWR.t26 28.5655
R2726 VPWR.n387 VPWR.t201 28.5655
R2727 VPWR.n387 VPWR.t203 28.5655
R2728 VPWR.n389 VPWR.t189 28.5655
R2729 VPWR.n389 VPWR.t197 28.5655
R2730 VPWR.n382 VPWR.t195 28.5655
R2731 VPWR.n382 VPWR.t193 28.5655
R2732 VPWR.n384 VPWR.t199 28.5655
R2733 VPWR.n384 VPWR.t187 28.5655
R2734 VPWR.n394 VPWR.t205 28.5655
R2735 VPWR.n394 VPWR.t191 28.5655
R2736 VPWR.n630 VPWR.t122 28.5655
R2737 VPWR.n630 VPWR.t126 28.5655
R2738 VPWR.n632 VPWR.t116 28.5655
R2739 VPWR.n632 VPWR.t114 28.5655
R2740 VPWR.n625 VPWR.t130 28.5655
R2741 VPWR.n625 VPWR.t120 28.5655
R2742 VPWR.n627 VPWR.t118 28.5655
R2743 VPWR.n627 VPWR.t124 28.5655
R2744 VPWR.n637 VPWR.t128 28.5655
R2745 VPWR.n637 VPWR.t132 28.5655
R2746 VPWR.n549 VPWR.t172 28.5655
R2747 VPWR.n549 VPWR.t176 28.5655
R2748 VPWR.n551 VPWR.t166 28.5655
R2749 VPWR.n551 VPWR.t184 28.5655
R2750 VPWR.n544 VPWR.t182 28.5655
R2751 VPWR.n544 VPWR.t168 28.5655
R2752 VPWR.n546 VPWR.t170 28.5655
R2753 VPWR.n546 VPWR.t174 28.5655
R2754 VPWR.n556 VPWR.t180 28.5655
R2755 VPWR.n556 VPWR.t178 28.5655
R2756 VPWR.n211 VPWR.t102 26.5955
R2757 VPWR.n211 VPWR.t99 26.5955
R2758 VPWR.n200 VPWR.t80 26.5955
R2759 VPWR.n200 VPWR.t33 26.5955
R2760 VPWR.n201 VPWR.t100 26.5955
R2761 VPWR.n201 VPWR.t34 26.5955
R2762 VPWR.n290 VPWR.t157 26.5955
R2763 VPWR.n290 VPWR.t159 26.5955
R2764 VPWR.n279 VPWR.t160 26.5955
R2765 VPWR.n279 VPWR.t96 26.5955
R2766 VPWR.n280 VPWR.t36 26.5955
R2767 VPWR.n280 VPWR.t37 26.5955
R2768 VPWR.n130 VPWR.t89 26.5955
R2769 VPWR.n130 VPWR.t49 26.5955
R2770 VPWR.n119 VPWR.t103 26.5955
R2771 VPWR.n119 VPWR.t228 26.5955
R2772 VPWR.n120 VPWR.t50 26.5955
R2773 VPWR.n120 VPWR.t87 26.5955
R2774 VPWR.n51 VPWR.t109 26.5955
R2775 VPWR.n51 VPWR.t10 26.5955
R2776 VPWR.n40 VPWR.t47 26.5955
R2777 VPWR.n40 VPWR.t11 26.5955
R2778 VPWR.n41 VPWR.t12 26.5955
R2779 VPWR.n41 VPWR.t110 26.5955
R2780 VPWR.n428 VPWR.t7 26.5955
R2781 VPWR.n428 VPWR.t9 26.5955
R2782 VPWR.n417 VPWR.t6 26.5955
R2783 VPWR.n417 VPWR.t4 26.5955
R2784 VPWR.n418 VPWR.t3 26.5955
R2785 VPWR.n418 VPWR.t1 26.5955
R2786 VPWR.n347 VPWR.t185 26.5955
R2787 VPWR.n347 VPWR.t288 26.5955
R2788 VPWR.n336 VPWR.t290 26.5955
R2789 VPWR.n336 VPWR.t133 26.5955
R2790 VPWR.n337 VPWR.t112 26.5955
R2791 VPWR.n337 VPWR.t135 26.5955
R2792 VPWR.n590 VPWR.t281 26.5955
R2793 VPWR.n590 VPWR.t283 26.5955
R2794 VPWR.n579 VPWR.t45 26.5955
R2795 VPWR.n579 VPWR.t43 26.5955
R2796 VPWR.n580 VPWR.t42 26.5955
R2797 VPWR.n580 VPWR.t44 26.5955
R2798 VPWR.n509 VPWR.t92 26.5955
R2799 VPWR.n509 VPWR.t83 26.5955
R2800 VPWR.n498 VPWR.t94 26.5955
R2801 VPWR.n498 VPWR.t84 26.5955
R2802 VPWR.n499 VPWR.t85 26.5955
R2803 VPWR.n499 VPWR.t93 26.5955
R2804 VPWR.n219 VPWR.n218 25.977
R2805 VPWR.n298 VPWR.n297 25.977
R2806 VPWR.n138 VPWR.n137 25.977
R2807 VPWR.n59 VPWR.n58 25.977
R2808 VPWR.n436 VPWR.n435 25.977
R2809 VPWR.n355 VPWR.n354 25.977
R2810 VPWR.n598 VPWR.n597 25.977
R2811 VPWR.n517 VPWR.n516 25.977
R2812 VPWR.n226 VPWR.n224 20.5561
R2813 VPWR.n233 VPWR.n231 20.5561
R2814 VPWR.n305 VPWR.n303 20.5561
R2815 VPWR.n312 VPWR.n310 20.5561
R2816 VPWR.n66 VPWR.n64 20.5561
R2817 VPWR.n73 VPWR.n71 20.5561
R2818 VPWR.n145 VPWR.n143 20.5561
R2819 VPWR.n152 VPWR.n150 20.5561
R2820 VPWR.n402 VPWR.n400 20.5561
R2821 VPWR.n409 VPWR.n407 20.5561
R2822 VPWR.n322 VPWR.n320 20.5561
R2823 VPWR.n329 VPWR.n327 20.5561
R2824 VPWR.n564 VPWR.n562 20.5561
R2825 VPWR.n571 VPWR.n569 20.5561
R2826 VPWR.n484 VPWR.n482 20.5561
R2827 VPWR.n491 VPWR.n489 20.5561
R2828 VPWR.n203 VPWR.n202 18.824
R2829 VPWR.n282 VPWR.n281 18.824
R2830 VPWR.n122 VPWR.n121 18.824
R2831 VPWR.n43 VPWR.n42 18.824
R2832 VPWR.n420 VPWR.n419 18.824
R2833 VPWR.n339 VPWR.n338 18.824
R2834 VPWR.n582 VPWR.n581 18.824
R2835 VPWR.n501 VPWR.n500 18.824
R2836 VPWR.n224 VPWR.n223 18.7435
R2837 VPWR.n231 VPWR.n230 18.7435
R2838 VPWR.n303 VPWR.n302 18.7435
R2839 VPWR.n310 VPWR.n309 18.7435
R2840 VPWR.n64 VPWR.n63 18.7435
R2841 VPWR.n71 VPWR.n70 18.7435
R2842 VPWR.n143 VPWR.n142 18.7435
R2843 VPWR.n150 VPWR.n149 18.7435
R2844 VPWR.n400 VPWR.n399 18.7435
R2845 VPWR.n407 VPWR.n406 18.7435
R2846 VPWR.n320 VPWR.n319 18.7435
R2847 VPWR.n327 VPWR.n326 18.7435
R2848 VPWR.n562 VPWR.n561 18.7435
R2849 VPWR.n569 VPWR.n568 18.7435
R2850 VPWR.n482 VPWR.n481 18.7435
R2851 VPWR.n489 VPWR.n488 18.7435
R2852 VPWR.n213 VPWR.n212 13.5534
R2853 VPWR.n292 VPWR.n291 13.5534
R2854 VPWR.n132 VPWR.n131 13.5534
R2855 VPWR.n53 VPWR.n52 13.5534
R2856 VPWR.n430 VPWR.n429 13.5534
R2857 VPWR.n349 VPWR.n348 13.5534
R2858 VPWR.n592 VPWR.n591 13.5534
R2859 VPWR.n511 VPWR.n510 13.5534
R2860 VPWR VPWR.n228 11.4981
R2861 VPWR VPWR.n235 11.4981
R2862 VPWR VPWR.n307 11.4981
R2863 VPWR VPWR.n314 11.4981
R2864 VPWR VPWR.n68 11.4981
R2865 VPWR VPWR.n75 11.4981
R2866 VPWR VPWR.n147 11.4981
R2867 VPWR VPWR.n154 11.4981
R2868 VPWR VPWR.n404 11.4981
R2869 VPWR VPWR.n411 11.4981
R2870 VPWR VPWR.n324 11.4981
R2871 VPWR VPWR.n331 11.4981
R2872 VPWR VPWR.n566 11.4981
R2873 VPWR VPWR.n573 11.4981
R2874 VPWR VPWR.n486 11.4981
R2875 VPWR VPWR.n493 11.4981
R2876 VPWR.n214 VPWR.n213 11.1829
R2877 VPWR.n293 VPWR.n292 11.1829
R2878 VPWR.n133 VPWR.n132 11.1829
R2879 VPWR.n54 VPWR.n53 11.1829
R2880 VPWR.n431 VPWR.n430 11.1829
R2881 VPWR.n350 VPWR.n349 11.1829
R2882 VPWR.n593 VPWR.n592 11.1829
R2883 VPWR.n512 VPWR.n511 11.1829
R2884 VPWR.n204 VPWR.n203 9.3005
R2885 VPWR.n205 VPWR.n202 9.3005
R2886 VPWR.n207 VPWR.n206 9.3005
R2887 VPWR.n209 VPWR.n198 9.3005
R2888 VPWR.n221 VPWR.n220 9.3005
R2889 VPWR.n219 VPWR.n199 9.3005
R2890 VPWR.n217 VPWR.n216 9.3005
R2891 VPWR.n215 VPWR.n212 9.3005
R2892 VPWR.n283 VPWR.n282 9.3005
R2893 VPWR.n284 VPWR.n281 9.3005
R2894 VPWR.n286 VPWR.n285 9.3005
R2895 VPWR.n288 VPWR.n277 9.3005
R2896 VPWR.n300 VPWR.n299 9.3005
R2897 VPWR.n298 VPWR.n278 9.3005
R2898 VPWR.n296 VPWR.n295 9.3005
R2899 VPWR.n294 VPWR.n291 9.3005
R2900 VPWR.n123 VPWR.n122 9.3005
R2901 VPWR.n124 VPWR.n121 9.3005
R2902 VPWR.n126 VPWR.n125 9.3005
R2903 VPWR.n128 VPWR.n117 9.3005
R2904 VPWR.n140 VPWR.n139 9.3005
R2905 VPWR.n138 VPWR.n118 9.3005
R2906 VPWR.n136 VPWR.n135 9.3005
R2907 VPWR.n134 VPWR.n131 9.3005
R2908 VPWR.n44 VPWR.n43 9.3005
R2909 VPWR.n45 VPWR.n42 9.3005
R2910 VPWR.n47 VPWR.n46 9.3005
R2911 VPWR.n49 VPWR.n38 9.3005
R2912 VPWR.n61 VPWR.n60 9.3005
R2913 VPWR.n59 VPWR.n39 9.3005
R2914 VPWR.n57 VPWR.n56 9.3005
R2915 VPWR.n55 VPWR.n52 9.3005
R2916 VPWR.n421 VPWR.n420 9.3005
R2917 VPWR.n422 VPWR.n419 9.3005
R2918 VPWR.n424 VPWR.n423 9.3005
R2919 VPWR.n426 VPWR.n415 9.3005
R2920 VPWR.n438 VPWR.n437 9.3005
R2921 VPWR.n436 VPWR.n416 9.3005
R2922 VPWR.n434 VPWR.n433 9.3005
R2923 VPWR.n432 VPWR.n429 9.3005
R2924 VPWR.n340 VPWR.n339 9.3005
R2925 VPWR.n341 VPWR.n338 9.3005
R2926 VPWR.n343 VPWR.n342 9.3005
R2927 VPWR.n345 VPWR.n334 9.3005
R2928 VPWR.n357 VPWR.n356 9.3005
R2929 VPWR.n355 VPWR.n335 9.3005
R2930 VPWR.n353 VPWR.n352 9.3005
R2931 VPWR.n351 VPWR.n348 9.3005
R2932 VPWR.n583 VPWR.n582 9.3005
R2933 VPWR.n584 VPWR.n581 9.3005
R2934 VPWR.n586 VPWR.n585 9.3005
R2935 VPWR.n588 VPWR.n577 9.3005
R2936 VPWR.n600 VPWR.n599 9.3005
R2937 VPWR.n598 VPWR.n578 9.3005
R2938 VPWR.n596 VPWR.n595 9.3005
R2939 VPWR.n594 VPWR.n591 9.3005
R2940 VPWR.n502 VPWR.n501 9.3005
R2941 VPWR.n503 VPWR.n500 9.3005
R2942 VPWR.n505 VPWR.n504 9.3005
R2943 VPWR.n507 VPWR.n496 9.3005
R2944 VPWR.n519 VPWR.n518 9.3005
R2945 VPWR.n517 VPWR.n497 9.3005
R2946 VPWR.n515 VPWR.n514 9.3005
R2947 VPWR.n513 VPWR.n510 9.3005
R2948 VPWR.n218 VPWR.n217 8.65932
R2949 VPWR.n297 VPWR.n296 8.65932
R2950 VPWR.n137 VPWR.n136 8.65932
R2951 VPWR.n58 VPWR.n57 8.65932
R2952 VPWR.n435 VPWR.n434 8.65932
R2953 VPWR.n354 VPWR.n353 8.65932
R2954 VPWR.n597 VPWR.n596 8.65932
R2955 VPWR.n516 VPWR.n515 8.65932
R2956 VPWR.n78 VPWR 5.89271
R2957 VPWR.n168 VPWR.n165 5.0005
R2958 VPWR.n174 VPWR.n165 5.0005
R2959 VPWR.n247 VPWR.n244 5.0005
R2960 VPWR.n253 VPWR.n244 5.0005
R2961 VPWR.n87 VPWR.n84 5.0005
R2962 VPWR.n93 VPWR.n84 5.0005
R2963 VPWR.n8 VPWR.n5 5.0005
R2964 VPWR.n14 VPWR.n5 5.0005
R2965 VPWR.n449 VPWR.n446 5.0005
R2966 VPWR.n455 VPWR.n446 5.0005
R2967 VPWR.n368 VPWR.n365 5.0005
R2968 VPWR.n374 VPWR.n365 5.0005
R2969 VPWR.n611 VPWR.n608 5.0005
R2970 VPWR.n617 VPWR.n608 5.0005
R2971 VPWR.n530 VPWR.n527 5.0005
R2972 VPWR.n536 VPWR.n527 5.0005
R2973 VPWR.n159 VPWR 4.95117
R2974 VPWR.n167 VPWR.n164 4.86892
R2975 VPWR.n166 VPWR.n164 4.86892
R2976 VPWR.n246 VPWR.n243 4.86892
R2977 VPWR.n245 VPWR.n243 4.86892
R2978 VPWR.n86 VPWR.n83 4.86892
R2979 VPWR.n85 VPWR.n83 4.86892
R2980 VPWR.n7 VPWR.n4 4.86892
R2981 VPWR.n6 VPWR.n4 4.86892
R2982 VPWR.n448 VPWR.n445 4.86892
R2983 VPWR.n447 VPWR.n445 4.86892
R2984 VPWR.n367 VPWR.n364 4.86892
R2985 VPWR.n366 VPWR.n364 4.86892
R2986 VPWR.n610 VPWR.n607 4.86892
R2987 VPWR.n609 VPWR.n607 4.86892
R2988 VPWR.n529 VPWR.n526 4.86892
R2989 VPWR.n528 VPWR.n526 4.86892
R2990 VPWR.n480 VPWR 3.8545
R2991 VPWR.n208 VPWR.n207 3.38874
R2992 VPWR.n287 VPWR.n286 3.38874
R2993 VPWR.n127 VPWR.n126 3.38874
R2994 VPWR.n48 VPWR.n47 3.38874
R2995 VPWR.n425 VPWR.n424 3.38874
R2996 VPWR.n344 VPWR.n343 3.38874
R2997 VPWR.n587 VPWR.n586 3.38874
R2998 VPWR.n506 VPWR.n505 3.38874
R2999 VPWR.n237 VPWR.n236 3.28283
R3000 VPWR.n316 VPWR.n315 3.28283
R3001 VPWR.n77 VPWR.n76 3.28283
R3002 VPWR.n156 VPWR.n155 3.28283
R3003 VPWR.n413 VPWR.n412 3.28283
R3004 VPWR.n333 VPWR.n332 3.28283
R3005 VPWR.n575 VPWR.n574 3.28283
R3006 VPWR.n495 VPWR.n494 3.28283
R3007 VPWR.n237 VPWR.n229 3.19667
R3008 VPWR.n316 VPWR.n308 3.19667
R3009 VPWR.n77 VPWR.n69 3.19667
R3010 VPWR.n156 VPWR.n148 3.19667
R3011 VPWR.n413 VPWR.n405 3.19667
R3012 VPWR.n333 VPWR.n325 3.19667
R3013 VPWR.n575 VPWR.n567 3.19667
R3014 VPWR.n495 VPWR.n487 3.19667
R3015 VPWR.n642 VPWR 2.7265
R3016 VPWR.n220 VPWR.n210 2.63579
R3017 VPWR.n299 VPWR.n289 2.63579
R3018 VPWR.n139 VPWR.n129 2.63579
R3019 VPWR.n60 VPWR.n50 2.63579
R3020 VPWR.n437 VPWR.n427 2.63579
R3021 VPWR.n356 VPWR.n346 2.63579
R3022 VPWR.n599 VPWR.n589 2.63579
R3023 VPWR.n518 VPWR.n508 2.63579
R3024 VPWR.n642 VPWR 2.5385
R3025 VPWR.n179 VPWR.n161 2.4755
R3026 VPWR.n169 VPWR.n161 2.4755
R3027 VPWR.n258 VPWR.n240 2.4755
R3028 VPWR.n248 VPWR.n240 2.4755
R3029 VPWR.n98 VPWR.n80 2.4755
R3030 VPWR.n88 VPWR.n80 2.4755
R3031 VPWR.n19 VPWR.n1 2.4755
R3032 VPWR.n9 VPWR.n1 2.4755
R3033 VPWR.n460 VPWR.n442 2.4755
R3034 VPWR.n450 VPWR.n442 2.4755
R3035 VPWR.n379 VPWR.n361 2.4755
R3036 VPWR.n369 VPWR.n361 2.4755
R3037 VPWR.n622 VPWR.n604 2.4755
R3038 VPWR.n612 VPWR.n604 2.4755
R3039 VPWR.n541 VPWR.n523 2.4755
R3040 VPWR.n531 VPWR.n523 2.4755
R3041 VPWR.n169 VPWR.n160 2.463
R3042 VPWR.n248 VPWR.n239 2.463
R3043 VPWR.n88 VPWR.n79 2.463
R3044 VPWR.n9 VPWR.n0 2.463
R3045 VPWR.n450 VPWR.n441 2.463
R3046 VPWR.n369 VPWR.n360 2.463
R3047 VPWR.n612 VPWR.n603 2.463
R3048 VPWR.n531 VPWR.n522 2.463
R3049 VPWR.n177 VPWR.n176 2.34227
R3050 VPWR.n176 VPWR.n175 2.34227
R3051 VPWR.n172 VPWR.n171 2.34227
R3052 VPWR.n173 VPWR.n172 2.34227
R3053 VPWR.n256 VPWR.n255 2.34227
R3054 VPWR.n255 VPWR.n254 2.34227
R3055 VPWR.n251 VPWR.n250 2.34227
R3056 VPWR.n252 VPWR.n251 2.34227
R3057 VPWR.n96 VPWR.n95 2.34227
R3058 VPWR.n95 VPWR.n94 2.34227
R3059 VPWR.n91 VPWR.n90 2.34227
R3060 VPWR.n92 VPWR.n91 2.34227
R3061 VPWR.n17 VPWR.n16 2.34227
R3062 VPWR.n16 VPWR.n15 2.34227
R3063 VPWR.n12 VPWR.n11 2.34227
R3064 VPWR.n13 VPWR.n12 2.34227
R3065 VPWR.n458 VPWR.n457 2.34227
R3066 VPWR.n457 VPWR.n456 2.34227
R3067 VPWR.n453 VPWR.n452 2.34227
R3068 VPWR.n454 VPWR.n453 2.34227
R3069 VPWR.n377 VPWR.n376 2.34227
R3070 VPWR.n376 VPWR.n375 2.34227
R3071 VPWR.n372 VPWR.n371 2.34227
R3072 VPWR.n373 VPWR.n372 2.34227
R3073 VPWR.n620 VPWR.n619 2.34227
R3074 VPWR.n619 VPWR.n618 2.34227
R3075 VPWR.n615 VPWR.n614 2.34227
R3076 VPWR.n616 VPWR.n615 2.34227
R3077 VPWR.n539 VPWR.n538 2.34227
R3078 VPWR.n538 VPWR.n537 2.34227
R3079 VPWR.n534 VPWR.n533 2.34227
R3080 VPWR.n535 VPWR.n534 2.34227
R3081 VPWR.n180 VPWR.n160 2.10363
R3082 VPWR.n259 VPWR.n239 2.10363
R3083 VPWR.n99 VPWR.n79 2.10363
R3084 VPWR.n20 VPWR.n0 2.10363
R3085 VPWR.n461 VPWR.n441 2.10363
R3086 VPWR.n380 VPWR.n360 2.10363
R3087 VPWR.n623 VPWR.n603 2.10363
R3088 VPWR.n542 VPWR.n522 2.10363
R3089 VPWR.n178 VPWR.n177 1.93989
R3090 VPWR.n257 VPWR.n256 1.93989
R3091 VPWR.n97 VPWR.n96 1.93989
R3092 VPWR.n18 VPWR.n17 1.93989
R3093 VPWR.n459 VPWR.n458 1.93989
R3094 VPWR.n378 VPWR.n377 1.93989
R3095 VPWR.n621 VPWR.n620 1.93989
R3096 VPWR.n540 VPWR.n539 1.93989
R3097 VPWR.n238 VPWR.n222 1.02714
R3098 VPWR.n317 VPWR.n301 1.02714
R3099 VPWR.n157 VPWR.n141 1.02714
R3100 VPWR.n78 VPWR.n62 1.02714
R3101 VPWR.n440 VPWR.n439 1.02714
R3102 VPWR.n359 VPWR.n358 1.02714
R3103 VPWR.n602 VPWR.n601 1.02714
R3104 VPWR.n521 VPWR.n520 1.02714
R3105 VPWR.n167 VPWR.n162 0.970197
R3106 VPWR.n171 VPWR.n170 0.970197
R3107 VPWR.n168 VPWR.n163 0.970197
R3108 VPWR.n246 VPWR.n241 0.970197
R3109 VPWR.n250 VPWR.n249 0.970197
R3110 VPWR.n247 VPWR.n242 0.970197
R3111 VPWR.n86 VPWR.n81 0.970197
R3112 VPWR.n90 VPWR.n89 0.970197
R3113 VPWR.n87 VPWR.n82 0.970197
R3114 VPWR.n7 VPWR.n2 0.970197
R3115 VPWR.n11 VPWR.n10 0.970197
R3116 VPWR.n8 VPWR.n3 0.970197
R3117 VPWR.n448 VPWR.n443 0.970197
R3118 VPWR.n452 VPWR.n451 0.970197
R3119 VPWR.n449 VPWR.n444 0.970197
R3120 VPWR.n367 VPWR.n362 0.970197
R3121 VPWR.n371 VPWR.n370 0.970197
R3122 VPWR.n368 VPWR.n363 0.970197
R3123 VPWR.n610 VPWR.n605 0.970197
R3124 VPWR.n614 VPWR.n613 0.970197
R3125 VPWR.n611 VPWR.n606 0.970197
R3126 VPWR.n529 VPWR.n524 0.970197
R3127 VPWR.n533 VPWR.n532 0.970197
R3128 VPWR.n530 VPWR.n525 0.970197
R3129 VPWR.n183 VPWR.n181 0.890989
R3130 VPWR.n262 VPWR.n260 0.890989
R3131 VPWR.n102 VPWR.n100 0.890989
R3132 VPWR.n23 VPWR.n21 0.890989
R3133 VPWR.n464 VPWR.n462 0.890989
R3134 VPWR.n383 VPWR.n381 0.890989
R3135 VPWR.n626 VPWR.n624 0.890989
R3136 VPWR.n545 VPWR.n543 0.890989
R3137 VPWR.n642 VPWR.n480 0.877833
R3138 VPWR.n480 VPWR.n318 0.8465
R3139 VPWR.n188 VPWR.n186 0.760446
R3140 VPWR.n267 VPWR.n265 0.760446
R3141 VPWR.n107 VPWR.n105 0.760446
R3142 VPWR.n28 VPWR.n26 0.760446
R3143 VPWR.n469 VPWR.n467 0.760446
R3144 VPWR.n388 VPWR.n386 0.760446
R3145 VPWR.n631 VPWR.n629 0.760446
R3146 VPWR.n550 VPWR.n548 0.760446
R3147 VPWR.n159 VPWR.n158 0.689833
R3148 VPWR.n190 VPWR.n188 0.40675
R3149 VPWR.n185 VPWR.n183 0.40675
R3150 VPWR.n195 VPWR.n185 0.40675
R3151 VPWR.n269 VPWR.n267 0.40675
R3152 VPWR.n264 VPWR.n262 0.40675
R3153 VPWR.n274 VPWR.n264 0.40675
R3154 VPWR.n109 VPWR.n107 0.40675
R3155 VPWR.n104 VPWR.n102 0.40675
R3156 VPWR.n114 VPWR.n104 0.40675
R3157 VPWR.n30 VPWR.n28 0.40675
R3158 VPWR.n25 VPWR.n23 0.40675
R3159 VPWR.n35 VPWR.n25 0.40675
R3160 VPWR.n471 VPWR.n469 0.40675
R3161 VPWR.n466 VPWR.n464 0.40675
R3162 VPWR.n476 VPWR.n466 0.40675
R3163 VPWR.n390 VPWR.n388 0.40675
R3164 VPWR.n385 VPWR.n383 0.40675
R3165 VPWR.n395 VPWR.n385 0.40675
R3166 VPWR.n633 VPWR.n631 0.40675
R3167 VPWR.n628 VPWR.n626 0.40675
R3168 VPWR.n638 VPWR.n628 0.40675
R3169 VPWR.n552 VPWR.n550 0.40675
R3170 VPWR.n547 VPWR.n545 0.40675
R3171 VPWR.n557 VPWR.n547 0.40675
R3172 VPWR.n521 VPWR.n495 0.397508
R3173 VPWR.n359 VPWR.n333 0.383506
R3174 VPWR.n180 VPWR.n179 0.359875
R3175 VPWR.n259 VPWR.n258 0.359875
R3176 VPWR.n99 VPWR.n98 0.359875
R3177 VPWR.n20 VPWR.n19 0.359875
R3178 VPWR.n461 VPWR.n460 0.359875
R3179 VPWR.n380 VPWR.n379 0.359875
R3180 VPWR.n623 VPWR.n622 0.359875
R3181 VPWR.n542 VPWR.n541 0.359875
R3182 VPWR.n157 VPWR.n156 0.3415
R3183 VPWR.n78 VPWR.n77 0.3415
R3184 VPWR.n317 VPWR.n316 0.3415
R3185 VPWR.n238 VPWR.n237 0.3415
R3186 VPWR.n414 VPWR.n413 0.3415
R3187 VPWR.n576 VPWR.n575 0.3415
R3188 VPWR.n163 VPWR.n161 0.258833
R3189 VPWR.n162 VPWR.n160 0.258833
R3190 VPWR.n242 VPWR.n240 0.258833
R3191 VPWR.n241 VPWR.n239 0.258833
R3192 VPWR.n82 VPWR.n80 0.258833
R3193 VPWR.n81 VPWR.n79 0.258833
R3194 VPWR.n3 VPWR.n1 0.258833
R3195 VPWR.n2 VPWR.n0 0.258833
R3196 VPWR.n444 VPWR.n442 0.258833
R3197 VPWR.n443 VPWR.n441 0.258833
R3198 VPWR.n363 VPWR.n361 0.258833
R3199 VPWR.n362 VPWR.n360 0.258833
R3200 VPWR.n606 VPWR.n604 0.258833
R3201 VPWR.n605 VPWR.n603 0.258833
R3202 VPWR.n525 VPWR.n523 0.258833
R3203 VPWR.n524 VPWR.n522 0.258833
R3204 VPWR.n195 VPWR.n193 0.208833
R3205 VPWR.n274 VPWR.n272 0.208833
R3206 VPWR.n114 VPWR.n112 0.208833
R3207 VPWR.n35 VPWR.n33 0.208833
R3208 VPWR.n476 VPWR.n474 0.208833
R3209 VPWR.n395 VPWR.n393 0.208833
R3210 VPWR.n638 VPWR.n636 0.208833
R3211 VPWR.n557 VPWR.n555 0.208833
R3212 VPWR.n193 VPWR.n190 0.188
R3213 VPWR.n272 VPWR.n269 0.188
R3214 VPWR.n112 VPWR.n109 0.188
R3215 VPWR.n33 VPWR.n30 0.188
R3216 VPWR.n474 VPWR.n471 0.188
R3217 VPWR.n393 VPWR.n390 0.188
R3218 VPWR.n636 VPWR.n633 0.188
R3219 VPWR.n555 VPWR.n552 0.188
R3220 VPWR.n193 VPWR.n192 0.1865
R3221 VPWR.n272 VPWR.n271 0.1865
R3222 VPWR.n112 VPWR.n111 0.1865
R3223 VPWR.n33 VPWR.n32 0.1865
R3224 VPWR.n474 VPWR.n473 0.1865
R3225 VPWR.n393 VPWR.n392 0.1865
R3226 VPWR.n636 VPWR.n635 0.1865
R3227 VPWR.n555 VPWR.n554 0.1865
R3228 VPWR.n560 VPWR.n521 0.184975
R3229 VPWR.n641 VPWR.n602 0.184975
R3230 VPWR.n642 VPWR 0.178395
R3231 VPWR.n576 VPWR 0.167428
R3232 VPWR.n398 VPWR.n359 0.138856
R3233 VPWR.n479 VPWR.n440 0.138856
R3234 VPWR.n480 VPWR 0.137564
R3235 VPWR.n170 VPWR.n169 0.121279
R3236 VPWR.n179 VPWR.n178 0.121279
R3237 VPWR.n249 VPWR.n248 0.121279
R3238 VPWR.n258 VPWR.n257 0.121279
R3239 VPWR.n89 VPWR.n88 0.121279
R3240 VPWR.n98 VPWR.n97 0.121279
R3241 VPWR.n10 VPWR.n9 0.121279
R3242 VPWR.n19 VPWR.n18 0.121279
R3243 VPWR.n451 VPWR.n450 0.121279
R3244 VPWR.n460 VPWR.n459 0.121279
R3245 VPWR.n370 VPWR.n369 0.121279
R3246 VPWR.n379 VPWR.n378 0.121279
R3247 VPWR.n613 VPWR.n612 0.121279
R3248 VPWR.n622 VPWR.n621 0.121279
R3249 VPWR.n532 VPWR.n531 0.121279
R3250 VPWR.n541 VPWR.n540 0.121279
R3251 VPWR.n205 VPWR.n204 0.120292
R3252 VPWR.n206 VPWR.n205 0.120292
R3253 VPWR.n206 VPWR.n198 0.120292
R3254 VPWR.n221 VPWR.n199 0.120292
R3255 VPWR.n216 VPWR.n199 0.120292
R3256 VPWR.n216 VPWR.n215 0.120292
R3257 VPWR.n215 VPWR.n214 0.120292
R3258 VPWR.n284 VPWR.n283 0.120292
R3259 VPWR.n285 VPWR.n284 0.120292
R3260 VPWR.n285 VPWR.n277 0.120292
R3261 VPWR.n300 VPWR.n278 0.120292
R3262 VPWR.n295 VPWR.n278 0.120292
R3263 VPWR.n295 VPWR.n294 0.120292
R3264 VPWR.n294 VPWR.n293 0.120292
R3265 VPWR.n124 VPWR.n123 0.120292
R3266 VPWR.n125 VPWR.n124 0.120292
R3267 VPWR.n125 VPWR.n117 0.120292
R3268 VPWR.n140 VPWR.n118 0.120292
R3269 VPWR.n135 VPWR.n118 0.120292
R3270 VPWR.n135 VPWR.n134 0.120292
R3271 VPWR.n134 VPWR.n133 0.120292
R3272 VPWR.n45 VPWR.n44 0.120292
R3273 VPWR.n46 VPWR.n45 0.120292
R3274 VPWR.n46 VPWR.n38 0.120292
R3275 VPWR.n61 VPWR.n39 0.120292
R3276 VPWR.n56 VPWR.n39 0.120292
R3277 VPWR.n56 VPWR.n55 0.120292
R3278 VPWR.n55 VPWR.n54 0.120292
R3279 VPWR.n422 VPWR.n421 0.120292
R3280 VPWR.n423 VPWR.n422 0.120292
R3281 VPWR.n423 VPWR.n415 0.120292
R3282 VPWR.n438 VPWR.n416 0.120292
R3283 VPWR.n433 VPWR.n416 0.120292
R3284 VPWR.n433 VPWR.n432 0.120292
R3285 VPWR.n432 VPWR.n431 0.120292
R3286 VPWR.n341 VPWR.n340 0.120292
R3287 VPWR.n342 VPWR.n341 0.120292
R3288 VPWR.n342 VPWR.n334 0.120292
R3289 VPWR.n357 VPWR.n335 0.120292
R3290 VPWR.n352 VPWR.n335 0.120292
R3291 VPWR.n352 VPWR.n351 0.120292
R3292 VPWR.n351 VPWR.n350 0.120292
R3293 VPWR.n584 VPWR.n583 0.120292
R3294 VPWR.n585 VPWR.n584 0.120292
R3295 VPWR.n585 VPWR.n577 0.120292
R3296 VPWR.n600 VPWR.n578 0.120292
R3297 VPWR.n595 VPWR.n578 0.120292
R3298 VPWR.n595 VPWR.n594 0.120292
R3299 VPWR.n594 VPWR.n593 0.120292
R3300 VPWR.n503 VPWR.n502 0.120292
R3301 VPWR.n504 VPWR.n503 0.120292
R3302 VPWR.n504 VPWR.n496 0.120292
R3303 VPWR.n519 VPWR.n497 0.120292
R3304 VPWR.n514 VPWR.n497 0.120292
R3305 VPWR.n514 VPWR.n513 0.120292
R3306 VPWR.n513 VPWR.n512 0.120292
R3307 VPWR.n222 VPWR.n221 0.115083
R3308 VPWR.n301 VPWR.n300 0.115083
R3309 VPWR.n141 VPWR.n140 0.115083
R3310 VPWR.n62 VPWR.n61 0.115083
R3311 VPWR.n439 VPWR.n438 0.115083
R3312 VPWR.n358 VPWR.n357 0.115083
R3313 VPWR.n601 VPWR.n600 0.115083
R3314 VPWR.n520 VPWR.n519 0.115083
R3315 VPWR.n414 VPWR 0.111772
R3316 VPWR VPWR.n560 0.109383
R3317 VPWR VPWR.n641 0.109383
R3318 VPWR.n196 VPWR.n195 0.0948367
R3319 VPWR.n275 VPWR.n274 0.0948367
R3320 VPWR.n115 VPWR.n114 0.0948367
R3321 VPWR.n36 VPWR.n35 0.0948367
R3322 VPWR.n477 VPWR.n476 0.0948367
R3323 VPWR.n396 VPWR.n395 0.0948367
R3324 VPWR.n639 VPWR.n638 0.0948367
R3325 VPWR.n558 VPWR.n557 0.0948367
R3326 VPWR VPWR.n398 0.0821625
R3327 VPWR VPWR.n479 0.0821625
R3328 VPWR.n196 VPWR.n180 0.0691538
R3329 VPWR.n275 VPWR.n259 0.0691538
R3330 VPWR.n115 VPWR.n99 0.0691538
R3331 VPWR.n36 VPWR.n20 0.0691538
R3332 VPWR.n477 VPWR.n461 0.0691538
R3333 VPWR.n396 VPWR.n380 0.0691538
R3334 VPWR.n639 VPWR.n623 0.0691538
R3335 VPWR.n558 VPWR.n542 0.0691538
R3336 VPWR.n197 VPWR.n196 0.0614341
R3337 VPWR.n276 VPWR.n275 0.0614341
R3338 VPWR.n116 VPWR.n115 0.0614341
R3339 VPWR.n37 VPWR.n36 0.0614341
R3340 VPWR.n478 VPWR.n477 0.0614341
R3341 VPWR.n397 VPWR.n396 0.0614341
R3342 VPWR.n640 VPWR.n639 0.0614341
R3343 VPWR.n559 VPWR.n558 0.0614341
R3344 VPWR.n158 VPWR 0.0613633
R3345 VPWR.n204 VPWR 0.0603958
R3346 VPWR.n283 VPWR 0.0603958
R3347 VPWR.n123 VPWR 0.0603958
R3348 VPWR.n44 VPWR 0.0603958
R3349 VPWR.n421 VPWR 0.0603958
R3350 VPWR.n340 VPWR 0.0603958
R3351 VPWR.n583 VPWR 0.0603958
R3352 VPWR.n502 VPWR 0.0603958
R3353 VPWR.n602 VPWR.n576 0.0565083
R3354 VPWR.n197 VPWR 0.0562442
R3355 VPWR.n276 VPWR 0.0562442
R3356 VPWR.n116 VPWR 0.0562442
R3357 VPWR.n37 VPWR 0.0562442
R3358 VPWR.n478 VPWR 0.0562442
R3359 VPWR.n397 VPWR 0.0562442
R3360 VPWR.n640 VPWR 0.0562442
R3361 VPWR.n559 VPWR 0.0562442
R3362 VPWR.n318 VPWR 0.0512194
R3363 VPWR.n229 VPWR 0.0459545
R3364 VPWR.n236 VPWR 0.0459545
R3365 VPWR.n308 VPWR 0.0459545
R3366 VPWR.n315 VPWR 0.0459545
R3367 VPWR.n69 VPWR 0.0459545
R3368 VPWR.n76 VPWR 0.0459545
R3369 VPWR.n148 VPWR 0.0459545
R3370 VPWR.n155 VPWR 0.0459545
R3371 VPWR.n405 VPWR 0.0459545
R3372 VPWR.n412 VPWR 0.0459545
R3373 VPWR.n325 VPWR 0.0459545
R3374 VPWR.n332 VPWR 0.0459545
R3375 VPWR.n567 VPWR 0.0459545
R3376 VPWR.n574 VPWR 0.0459545
R3377 VPWR.n487 VPWR 0.0459545
R3378 VPWR.n494 VPWR 0.0459545
R3379 VPWR.n440 VPWR.n414 0.0425062
R3380 VPWR.n229 VPWR 0.0338333
R3381 VPWR.n236 VPWR 0.0338333
R3382 VPWR.n308 VPWR 0.0338333
R3383 VPWR.n315 VPWR 0.0338333
R3384 VPWR.n69 VPWR 0.0338333
R3385 VPWR.n76 VPWR 0.0338333
R3386 VPWR.n148 VPWR 0.0338333
R3387 VPWR.n155 VPWR 0.0338333
R3388 VPWR.n405 VPWR 0.0338333
R3389 VPWR.n412 VPWR 0.0338333
R3390 VPWR.n325 VPWR 0.0338333
R3391 VPWR.n332 VPWR 0.0338333
R3392 VPWR.n567 VPWR 0.0338333
R3393 VPWR.n574 VPWR 0.0338333
R3394 VPWR.n487 VPWR 0.0338333
R3395 VPWR.n494 VPWR 0.0338333
R3396 VPWR.n214 VPWR 0.0226354
R3397 VPWR.n293 VPWR 0.0226354
R3398 VPWR.n133 VPWR 0.0226354
R3399 VPWR.n54 VPWR 0.0226354
R3400 VPWR.n431 VPWR 0.0226354
R3401 VPWR.n350 VPWR 0.0226354
R3402 VPWR.n593 VPWR 0.0226354
R3403 VPWR.n512 VPWR 0.0226354
R3404 VPWR VPWR.n642 0.006375
R3405 VPWR.n78 VPWR.n37 0.00599114
R3406 VPWR.n157 VPWR.n116 0.00599114
R3407 VPWR.n317 VPWR.n276 0.00599114
R3408 VPWR.n238 VPWR.n197 0.00599114
R3409 VPWR.n398 VPWR.n397 0.00599114
R3410 VPWR.n479 VPWR.n478 0.00599114
R3411 VPWR.n560 VPWR.n559 0.00599114
R3412 VPWR.n641 VPWR.n640 0.00599114
R3413 VPWR.n222 VPWR.n198 0.00570833
R3414 VPWR.n301 VPWR.n277 0.00570833
R3415 VPWR.n141 VPWR.n117 0.00570833
R3416 VPWR.n62 VPWR.n38 0.00570833
R3417 VPWR.n439 VPWR.n415 0.00570833
R3418 VPWR.n358 VPWR.n334 0.00570833
R3419 VPWR.n601 VPWR.n577 0.00570833
R3420 VPWR.n520 VPWR.n496 0.00570833
R3421 VPWR.n480 VPWR 0.00490625
R3422 VPWR.n238 VPWR.n159 0.00211964
R3423 VPWR VPWR.n317 0.00099705
R3424 VPWR VPWR.n157 0.000926043
R3425 VPWR.n158 VPWR 0.000834748
R3426 VPWR.n318 VPWR 0.000831367
R3427 VPWR.n157 VPWR.n78 0.000699496
R3428 VPWR.n317 VPWR.n238 0.000628489
R3429 ui_in[6].n2 ui_in[6].t1 212.081
R3430 ui_in[6].n1 ui_in[6].t4 212.081
R3431 ui_in[6].n6 ui_in[6].t6 212.081
R3432 ui_in[6].n0 ui_in[6].t7 212.081
R3433 ui_in[6].n11 ui_in[6].t5 212.081
R3434 ui_in[6].n17 ui_in[6].t0 212.081
R3435 ui_in[6].n12 ui_in[6].t2 212.081
R3436 ui_in[6].n13 ui_in[6].t18 212.081
R3437 ui_in[6] ui_in[6].n14 163.264
R3438 ui_in[6].n16 ui_in[6].n15 152
R3439 ui_in[6].n19 ui_in[6].n18 152
R3440 ui_in[6].n10 ui_in[6].n9 152
R3441 ui_in[6].n8 ui_in[6].n7 152
R3442 ui_in[6].n5 ui_in[6].n4 152
R3443 ui_in[6] ui_in[6].n3 152
R3444 ui_in[6].n2 ui_in[6].t12 139.78
R3445 ui_in[6].n1 ui_in[6].t14 139.78
R3446 ui_in[6].n6 ui_in[6].t16 139.78
R3447 ui_in[6].n0 ui_in[6].t17 139.78
R3448 ui_in[6].n11 ui_in[6].t15 139.78
R3449 ui_in[6].n17 ui_in[6].t11 139.78
R3450 ui_in[6].n12 ui_in[6].t13 139.78
R3451 ui_in[6].n13 ui_in[6].t9 139.78
R3452 ui_in[6].n24 ui_in[6].t19 120.23
R3453 ui_in[6].n24 ui_in[6].t3 120.228
R3454 ui_in[6].n21 ui_in[6].t8 118.061
R3455 ui_in[6].n21 ui_in[6].t10 118.058
R3456 ui_in[6].n3 ui_in[6].n2 30.6732
R3457 ui_in[6].n3 ui_in[6].n1 30.6732
R3458 ui_in[6].n5 ui_in[6].n1 30.6732
R3459 ui_in[6].n6 ui_in[6].n5 30.6732
R3460 ui_in[6].n7 ui_in[6].n6 30.6732
R3461 ui_in[6].n7 ui_in[6].n0 30.6732
R3462 ui_in[6].n10 ui_in[6].n0 30.6732
R3463 ui_in[6].n11 ui_in[6].n10 30.6732
R3464 ui_in[6].n18 ui_in[6].n11 30.6732
R3465 ui_in[6].n18 ui_in[6].n17 30.6732
R3466 ui_in[6].n17 ui_in[6].n16 30.6732
R3467 ui_in[6].n16 ui_in[6].n12 30.6732
R3468 ui_in[6].n14 ui_in[6].n12 30.6732
R3469 ui_in[6].n14 ui_in[6].n13 30.6732
R3470 ui_in[6].n4 ui_in[6] 21.5045
R3471 ui_in[6].n8 ui_in[6] 19.4565
R3472 ui_in[6].n9 ui_in[6] 17.4085
R3473 ui_in[6].n15 ui_in[6] 13.3125
R3474 ui_in[6].n20 ui_in[6].n19 13.0565
R3475 ui_in[6].n15 ui_in[6] 10.2405
R3476 ui_in[6].n19 ui_in[6] 8.1925
R3477 ui_in[6].n9 ui_in[6] 6.1445
R3478 ui_in[6] ui_in[6].n8 4.0965
R3479 ui_in[6].n23 ui_in[6].n20 3.2054
R3480 ui_in[6].n20 ui_in[6] 2.3045
R3481 ui_in[6].n4 ui_in[6] 2.0485
R3482 ui_in[6].n22 ui_in[6].n21 0.528909
R3483 ui_in[6].n25 ui_in[6].n24 0.506182
R3484 ui_in[6].n26 ui_in[6].n25 0.42675
R3485 ui_in[6].n26 ui_in[6].n23 0.342556
R3486 ui_in[6].n23 ui_in[6].n22 0.3415
R3487 ui_in[6].n25 ui_in[6] 0.170955
R3488 ui_in[6].n22 ui_in[6] 0.148227
R3489 ui_in[6] ui_in[6].n26 0.01225
R3490 ui_in[3].n2 ui_in[3].t17 212.081
R3491 ui_in[3].n1 ui_in[3].t15 212.081
R3492 ui_in[3].n6 ui_in[3].t16 212.081
R3493 ui_in[3].n0 ui_in[3].t12 212.081
R3494 ui_in[3].n11 ui_in[3].t8 212.081
R3495 ui_in[3].n17 ui_in[3].t9 212.081
R3496 ui_in[3].n12 ui_in[3].t11 212.081
R3497 ui_in[3].n13 ui_in[3].t13 212.081
R3498 ui_in[3] ui_in[3].n14 163.264
R3499 ui_in[3].n16 ui_in[3].n15 152
R3500 ui_in[3].n19 ui_in[3].n18 152
R3501 ui_in[3].n10 ui_in[3].n9 152
R3502 ui_in[3].n8 ui_in[3].n7 152
R3503 ui_in[3].n5 ui_in[3].n4 152
R3504 ui_in[3] ui_in[3].n3 152
R3505 ui_in[3].n2 ui_in[3].t7 139.78
R3506 ui_in[3].n1 ui_in[3].t5 139.78
R3507 ui_in[3].n6 ui_in[3].t6 139.78
R3508 ui_in[3].n0 ui_in[3].t2 139.78
R3509 ui_in[3].n11 ui_in[3].t18 139.78
R3510 ui_in[3].n17 ui_in[3].t19 139.78
R3511 ui_in[3].n12 ui_in[3].t1 139.78
R3512 ui_in[3].n13 ui_in[3].t3 139.78
R3513 ui_in[3].n24 ui_in[3].t0 120.23
R3514 ui_in[3].n24 ui_in[3].t10 120.228
R3515 ui_in[3].n21 ui_in[3].t14 118.061
R3516 ui_in[3].n21 ui_in[3].t4 118.058
R3517 ui_in[3].n3 ui_in[3].n2 30.6732
R3518 ui_in[3].n3 ui_in[3].n1 30.6732
R3519 ui_in[3].n5 ui_in[3].n1 30.6732
R3520 ui_in[3].n6 ui_in[3].n5 30.6732
R3521 ui_in[3].n7 ui_in[3].n6 30.6732
R3522 ui_in[3].n7 ui_in[3].n0 30.6732
R3523 ui_in[3].n10 ui_in[3].n0 30.6732
R3524 ui_in[3].n11 ui_in[3].n10 30.6732
R3525 ui_in[3].n18 ui_in[3].n11 30.6732
R3526 ui_in[3].n18 ui_in[3].n17 30.6732
R3527 ui_in[3].n17 ui_in[3].n16 30.6732
R3528 ui_in[3].n16 ui_in[3].n12 30.6732
R3529 ui_in[3].n14 ui_in[3].n12 30.6732
R3530 ui_in[3].n14 ui_in[3].n13 30.6732
R3531 ui_in[3].n4 ui_in[3] 21.5045
R3532 ui_in[3].n8 ui_in[3] 19.4565
R3533 ui_in[3].n9 ui_in[3] 17.4085
R3534 ui_in[3].n15 ui_in[3] 13.3125
R3535 ui_in[3].n20 ui_in[3].n19 13.0565
R3536 ui_in[3].n15 ui_in[3] 10.2405
R3537 ui_in[3].n19 ui_in[3] 8.1925
R3538 ui_in[3].n9 ui_in[3] 6.1445
R3539 ui_in[3] ui_in[3].n8 4.0965
R3540 ui_in[3].n23 ui_in[3].n20 3.2054
R3541 ui_in[3].n20 ui_in[3] 2.3045
R3542 ui_in[3].n4 ui_in[3] 2.0485
R3543 ui_in[3].n22 ui_in[3].n21 0.528909
R3544 ui_in[3].n25 ui_in[3].n24 0.506182
R3545 ui_in[3].n26 ui_in[3].n25 0.42675
R3546 ui_in[3].n26 ui_in[3].n23 0.342556
R3547 ui_in[3].n23 ui_in[3].n22 0.3415
R3548 ui_in[3].n25 ui_in[3] 0.170955
R3549 ui_in[3].n22 ui_in[3] 0.148227
R3550 ui_in[3] ui_in[3].n26 0.01225
R3551 distortionUnit_5.IN.n0 distortionUnit_5.IN.t0 223.565
R3552 distortionUnit_5.IN.n3 distortionUnit_5.IN.t1 223.565
R3553 distortionUnit_5.IN.n14 distortionUnit_5.IN.n12 199.941
R3554 distortionUnit_5.IN.n8 distortionUnit_5.IN.n6 199.941
R3555 distortionUnit_5.IN.n19 distortionUnit_5.IN.t14 118.769
R3556 distortionUnit_5.IN.n22 distortionUnit_5.IN.t12 118.621
R3557 distortionUnit_5.IN.n21 distortionUnit_5.IN.t16 118.005
R3558 distortionUnit_5.IN.n20 distortionUnit_5.IN.t15 118.005
R3559 distortionUnit_5.IN.n19 distortionUnit_5.IN.t13 118.005
R3560 distortionUnit_5.IN.n2 distortionUnit_5.IN.n1 90.2112
R3561 distortionUnit_5.IN.n13 distortionUnit_5.IN.t8 83.7234
R3562 distortionUnit_5.IN.n15 distortionUnit_5.IN.t9 83.7234
R3563 distortionUnit_5.IN.n7 distortionUnit_5.IN.t7 83.7234
R3564 distortionUnit_5.IN.n9 distortionUnit_5.IN.t6 83.7234
R3565 distortionUnit_5.IN.n2 distortionUnit_5.IN.n0 66.2405
R3566 distortionUnit_5.IN.n3 distortionUnit_5.IN.n2 63.2157
R3567 distortionUnit_5.IN.n12 distortionUnit_5.IN.t5 28.5655
R3568 distortionUnit_5.IN.n12 distortionUnit_5.IN.t4 28.5655
R3569 distortionUnit_5.IN.n6 distortionUnit_5.IN.t11 28.5655
R3570 distortionUnit_5.IN.n6 distortionUnit_5.IN.t10 28.5655
R3571 distortionUnit_5.IN.n1 distortionUnit_5.IN.t2 17.4005
R3572 distortionUnit_5.IN.n1 distortionUnit_5.IN.t3 17.4005
R3573 distortionUnit_5.IN.n4 distortionUnit_5.IN.n0 5.54823
R3574 distortionUnit_5.IN.n4 distortionUnit_5.IN.n3 5.18686
R3575 distortionUnit_5.IN distortionUnit_5.IN.n18 4.9113
R3576 distortionUnit_5.IN distortionUnit_5.IN.n23 4.4438
R3577 distortionUnit_5.IN distortionUnit_5.IN.n22 2.77717
R3578 distortionUnit_5.IN.n20 distortionUnit_5.IN.n19 2.66195
R3579 distortionUnit_5.IN.n22 distortionUnit_5.IN.n21 1.71868
R3580 distortionUnit_5.IN.n17 distortionUnit_5.IN.n10 1.15259
R3581 distortionUnit_5.IN.n17 distortionUnit_5.IN.n16 0.938152
R3582 distortionUnit_5.IN.n21 distortionUnit_5.IN.n20 0.764886
R3583 distortionUnit_5.IN.n13 distortionUnit_5.IN.n11 0.5005
R3584 distortionUnit_5.IN.n16 distortionUnit_5.IN.n15 0.5005
R3585 distortionUnit_5.IN.n7 distortionUnit_5.IN.n5 0.5005
R3586 distortionUnit_5.IN.n10 distortionUnit_5.IN.n9 0.5005
R3587 distortionUnit_5.IN.n23 distortionUnit_5.IN 0.490406
R3588 distortionUnit_5.IN.n15 distortionUnit_5.IN.n14 0.478385
R3589 distortionUnit_5.IN.n14 distortionUnit_5.IN.n13 0.478385
R3590 distortionUnit_5.IN.n9 distortionUnit_5.IN.n8 0.478385
R3591 distortionUnit_5.IN.n8 distortionUnit_5.IN.n7 0.478385
R3592 distortionUnit_5.IN.n16 distortionUnit_5.IN.n11 0.364136
R3593 distortionUnit_5.IN.n10 distortionUnit_5.IN.n5 0.364136
R3594 distortionUnit_5.IN.n11 distortionUnit_5.IN 0.244818
R3595 distortionUnit_5.IN.n5 distortionUnit_5.IN 0.244818
R3596 distortionUnit_5.IN distortionUnit_5.IN.n4 0.244818
R3597 distortionUnit_5.IN.n18 distortionUnit_5.IN 0.150313
R3598 distortionUnit_5.IN.n18 distortionUnit_5.IN 0.024
R3599 distortionUnit_5.IN distortionUnit_5.IN.n17 0.0137188
R3600 distortionUnit_5.IN.n23 distortionUnit_5.IN 0.0129412
R3601 ui_in[7].n2 ui_in[7].t5 212.081
R3602 ui_in[7].n1 ui_in[7].t9 212.081
R3603 ui_in[7].n6 ui_in[7].t3 212.081
R3604 ui_in[7].n0 ui_in[7].t4 212.081
R3605 ui_in[7].n11 ui_in[7].t8 212.081
R3606 ui_in[7].n17 ui_in[7].t2 212.081
R3607 ui_in[7].n12 ui_in[7].t6 212.081
R3608 ui_in[7].n13 ui_in[7].t1 212.081
R3609 ui_in[7] ui_in[7].n14 163.264
R3610 ui_in[7].n16 ui_in[7].n15 152
R3611 ui_in[7].n19 ui_in[7].n18 152
R3612 ui_in[7].n10 ui_in[7].n9 152
R3613 ui_in[7].n8 ui_in[7].n7 152
R3614 ui_in[7].n5 ui_in[7].n4 152
R3615 ui_in[7] ui_in[7].n3 152
R3616 ui_in[7].n2 ui_in[7].t15 139.78
R3617 ui_in[7].n1 ui_in[7].t18 139.78
R3618 ui_in[7].n6 ui_in[7].t13 139.78
R3619 ui_in[7].n0 ui_in[7].t14 139.78
R3620 ui_in[7].n11 ui_in[7].t17 139.78
R3621 ui_in[7].n17 ui_in[7].t12 139.78
R3622 ui_in[7].n12 ui_in[7].t16 139.78
R3623 ui_in[7].n13 ui_in[7].t11 139.78
R3624 ui_in[7].n24 ui_in[7].t19 120.23
R3625 ui_in[7].n24 ui_in[7].t0 120.228
R3626 ui_in[7].n21 ui_in[7].t7 118.061
R3627 ui_in[7].n21 ui_in[7].t10 118.058
R3628 ui_in[7].n3 ui_in[7].n2 30.6732
R3629 ui_in[7].n3 ui_in[7].n1 30.6732
R3630 ui_in[7].n5 ui_in[7].n1 30.6732
R3631 ui_in[7].n6 ui_in[7].n5 30.6732
R3632 ui_in[7].n7 ui_in[7].n6 30.6732
R3633 ui_in[7].n7 ui_in[7].n0 30.6732
R3634 ui_in[7].n10 ui_in[7].n0 30.6732
R3635 ui_in[7].n11 ui_in[7].n10 30.6732
R3636 ui_in[7].n18 ui_in[7].n11 30.6732
R3637 ui_in[7].n18 ui_in[7].n17 30.6732
R3638 ui_in[7].n17 ui_in[7].n16 30.6732
R3639 ui_in[7].n16 ui_in[7].n12 30.6732
R3640 ui_in[7].n14 ui_in[7].n12 30.6732
R3641 ui_in[7].n14 ui_in[7].n13 30.6732
R3642 ui_in[7].n4 ui_in[7] 21.5045
R3643 ui_in[7].n8 ui_in[7] 19.4565
R3644 ui_in[7].n9 ui_in[7] 17.4085
R3645 ui_in[7].n15 ui_in[7] 13.3125
R3646 ui_in[7].n20 ui_in[7].n19 13.0565
R3647 ui_in[7].n15 ui_in[7] 10.2405
R3648 ui_in[7].n19 ui_in[7] 8.1925
R3649 ui_in[7].n9 ui_in[7] 6.1445
R3650 ui_in[7] ui_in[7].n8 4.0965
R3651 ui_in[7].n23 ui_in[7].n20 3.2054
R3652 ui_in[7].n20 ui_in[7] 2.3045
R3653 ui_in[7].n4 ui_in[7] 2.0485
R3654 ui_in[7].n22 ui_in[7].n21 0.528909
R3655 ui_in[7].n25 ui_in[7].n24 0.506182
R3656 ui_in[7].n26 ui_in[7].n25 0.42675
R3657 ui_in[7].n26 ui_in[7].n23 0.342556
R3658 ui_in[7].n23 ui_in[7].n22 0.3415
R3659 ui_in[7].n25 ui_in[7] 0.170955
R3660 ui_in[7].n22 ui_in[7] 0.148227
R3661 ui_in[7] ui_in[7].n26 0.01225
R3662 ua[1].n9 ua[1].n7 199.941
R3663 ua[1].n3 ua[1].n1 199.941
R3664 ua[1].n8 ua[1].t6 83.7234
R3665 ua[1].n10 ua[1].t7 83.7234
R3666 ua[1].n2 ua[1].t0 83.7234
R3667 ua[1].n4 ua[1].t1 83.7234
R3668 ua[1].n7 ua[1].t2 28.5655
R3669 ua[1].n7 ua[1].t3 28.5655
R3670 ua[1].n1 ua[1].t5 28.5655
R3671 ua[1].n1 ua[1].t4 28.5655
R3672 ua[1].n13 ua[1] 4.9995
R3673 ua[1].n12 ua[1].n5 1.15259
R3674 ua[1].n12 ua[1].n11 0.938152
R3675 ua[1].n8 ua[1].n6 0.5005
R3676 ua[1].n11 ua[1].n10 0.5005
R3677 ua[1].n2 ua[1].n0 0.5005
R3678 ua[1].n5 ua[1].n4 0.5005
R3679 ua[1].n10 ua[1].n9 0.478385
R3680 ua[1].n9 ua[1].n8 0.478385
R3681 ua[1].n4 ua[1].n3 0.478385
R3682 ua[1].n3 ua[1].n2 0.478385
R3683 ua[1].n11 ua[1].n6 0.364136
R3684 ua[1].n5 ua[1].n0 0.364136
R3685 ua[1].n6 ua[1] 0.244818
R3686 ua[1].n0 ua[1] 0.244818
R3687 ua[1].n13 ua[1] 0.150313
R3688 ua[1] ua[1].n13 0.024
R3689 ua[1] ua[1].n12 0.0137188
R3690 ui_in[0].n2 ui_in[0].t18 212.081
R3691 ui_in[0].n1 ui_in[0].t12 212.081
R3692 ui_in[0].n6 ui_in[0].t14 212.081
R3693 ui_in[0].n0 ui_in[0].t17 212.081
R3694 ui_in[0].n11 ui_in[0].t0 212.081
R3695 ui_in[0].n17 ui_in[0].t16 212.081
R3696 ui_in[0].n12 ui_in[0].t11 212.081
R3697 ui_in[0].n13 ui_in[0].t13 212.081
R3698 ui_in[0] ui_in[0].n14 163.264
R3699 ui_in[0].n16 ui_in[0].n15 152
R3700 ui_in[0].n19 ui_in[0].n18 152
R3701 ui_in[0].n10 ui_in[0].n9 152
R3702 ui_in[0].n8 ui_in[0].n7 152
R3703 ui_in[0].n5 ui_in[0].n4 152
R3704 ui_in[0] ui_in[0].n3 152
R3705 ui_in[0].n2 ui_in[0].t9 139.78
R3706 ui_in[0].n1 ui_in[0].t3 139.78
R3707 ui_in[0].n6 ui_in[0].t5 139.78
R3708 ui_in[0].n0 ui_in[0].t8 139.78
R3709 ui_in[0].n11 ui_in[0].t10 139.78
R3710 ui_in[0].n17 ui_in[0].t7 139.78
R3711 ui_in[0].n12 ui_in[0].t1 139.78
R3712 ui_in[0].n13 ui_in[0].t4 139.78
R3713 ui_in[0].n24 ui_in[0].t15 120.23
R3714 ui_in[0].n24 ui_in[0].t19 120.228
R3715 ui_in[0].n21 ui_in[0].t2 118.061
R3716 ui_in[0].n21 ui_in[0].t6 118.058
R3717 ui_in[0].n3 ui_in[0].n2 30.6732
R3718 ui_in[0].n3 ui_in[0].n1 30.6732
R3719 ui_in[0].n5 ui_in[0].n1 30.6732
R3720 ui_in[0].n6 ui_in[0].n5 30.6732
R3721 ui_in[0].n7 ui_in[0].n6 30.6732
R3722 ui_in[0].n7 ui_in[0].n0 30.6732
R3723 ui_in[0].n10 ui_in[0].n0 30.6732
R3724 ui_in[0].n11 ui_in[0].n10 30.6732
R3725 ui_in[0].n18 ui_in[0].n11 30.6732
R3726 ui_in[0].n18 ui_in[0].n17 30.6732
R3727 ui_in[0].n17 ui_in[0].n16 30.6732
R3728 ui_in[0].n16 ui_in[0].n12 30.6732
R3729 ui_in[0].n14 ui_in[0].n12 30.6732
R3730 ui_in[0].n14 ui_in[0].n13 30.6732
R3731 ui_in[0].n4 ui_in[0] 21.5045
R3732 ui_in[0].n8 ui_in[0] 19.4565
R3733 ui_in[0].n9 ui_in[0] 17.4085
R3734 ui_in[0].n15 ui_in[0] 13.3125
R3735 ui_in[0].n20 ui_in[0].n19 13.0565
R3736 ui_in[0].n15 ui_in[0] 10.2405
R3737 ui_in[0].n19 ui_in[0] 8.1925
R3738 ui_in[0].n9 ui_in[0] 6.1445
R3739 ui_in[0] ui_in[0].n8 4.0965
R3740 ui_in[0].n23 ui_in[0].n20 3.2054
R3741 ui_in[0].n20 ui_in[0] 2.3045
R3742 ui_in[0].n4 ui_in[0] 2.0485
R3743 ui_in[0].n22 ui_in[0].n21 0.528909
R3744 ui_in[0].n25 ui_in[0].n24 0.506182
R3745 ui_in[0].n26 ui_in[0].n25 0.42675
R3746 ui_in[0].n26 ui_in[0].n23 0.342556
R3747 ui_in[0].n23 ui_in[0].n22 0.3415
R3748 ui_in[0].n25 ui_in[0] 0.170955
R3749 ui_in[0].n22 ui_in[0] 0.148227
R3750 ui_in[0] ui_in[0].n26 0.01225
R3751 ui_in[2].n2 ui_in[2].t5 212.081
R3752 ui_in[2].n1 ui_in[2].t1 212.081
R3753 ui_in[2].n6 ui_in[2].t10 212.081
R3754 ui_in[2].n0 ui_in[2].t4 212.081
R3755 ui_in[2].n11 ui_in[2].t9 212.081
R3756 ui_in[2].n17 ui_in[2].t3 212.081
R3757 ui_in[2].n12 ui_in[2].t0 212.081
R3758 ui_in[2].n13 ui_in[2].t2 212.081
R3759 ui_in[2] ui_in[2].n14 163.264
R3760 ui_in[2].n16 ui_in[2].n15 152
R3761 ui_in[2].n19 ui_in[2].n18 152
R3762 ui_in[2].n10 ui_in[2].n9 152
R3763 ui_in[2].n8 ui_in[2].n7 152
R3764 ui_in[2].n5 ui_in[2].n4 152
R3765 ui_in[2] ui_in[2].n3 152
R3766 ui_in[2].n2 ui_in[2].t13 139.78
R3767 ui_in[2].n1 ui_in[2].t7 139.78
R3768 ui_in[2].n6 ui_in[2].t16 139.78
R3769 ui_in[2].n0 ui_in[2].t12 139.78
R3770 ui_in[2].n11 ui_in[2].t15 139.78
R3771 ui_in[2].n17 ui_in[2].t11 139.78
R3772 ui_in[2].n12 ui_in[2].t6 139.78
R3773 ui_in[2].n13 ui_in[2].t8 139.78
R3774 ui_in[2].n24 ui_in[2].t14 120.23
R3775 ui_in[2].n24 ui_in[2].t17 120.228
R3776 ui_in[2].n21 ui_in[2].t18 118.061
R3777 ui_in[2].n21 ui_in[2].t19 118.058
R3778 ui_in[2].n3 ui_in[2].n2 30.6732
R3779 ui_in[2].n3 ui_in[2].n1 30.6732
R3780 ui_in[2].n5 ui_in[2].n1 30.6732
R3781 ui_in[2].n6 ui_in[2].n5 30.6732
R3782 ui_in[2].n7 ui_in[2].n6 30.6732
R3783 ui_in[2].n7 ui_in[2].n0 30.6732
R3784 ui_in[2].n10 ui_in[2].n0 30.6732
R3785 ui_in[2].n11 ui_in[2].n10 30.6732
R3786 ui_in[2].n18 ui_in[2].n11 30.6732
R3787 ui_in[2].n18 ui_in[2].n17 30.6732
R3788 ui_in[2].n17 ui_in[2].n16 30.6732
R3789 ui_in[2].n16 ui_in[2].n12 30.6732
R3790 ui_in[2].n14 ui_in[2].n12 30.6732
R3791 ui_in[2].n14 ui_in[2].n13 30.6732
R3792 ui_in[2].n4 ui_in[2] 21.5045
R3793 ui_in[2].n8 ui_in[2] 19.4565
R3794 ui_in[2].n9 ui_in[2] 17.4085
R3795 ui_in[2].n15 ui_in[2] 13.3125
R3796 ui_in[2].n20 ui_in[2].n19 13.0565
R3797 ui_in[2].n15 ui_in[2] 10.2405
R3798 ui_in[2].n19 ui_in[2] 8.1925
R3799 ui_in[2].n9 ui_in[2] 6.1445
R3800 ui_in[2] ui_in[2].n8 4.0965
R3801 ui_in[2].n23 ui_in[2].n20 3.2054
R3802 ui_in[2].n20 ui_in[2] 2.3045
R3803 ui_in[2].n4 ui_in[2] 2.0485
R3804 ui_in[2].n22 ui_in[2].n21 0.528909
R3805 ui_in[2].n25 ui_in[2].n24 0.506182
R3806 ui_in[2].n26 ui_in[2].n25 0.42675
R3807 ui_in[2].n26 ui_in[2].n23 0.342556
R3808 ui_in[2].n23 ui_in[2].n22 0.3415
R3809 ui_in[2].n25 ui_in[2] 0.170955
R3810 ui_in[2].n22 ui_in[2] 0.148227
R3811 ui_in[2] ui_in[2].n26 0.01225
R3812 ui_in[5].n2 ui_in[5].t19 212.081
R3813 ui_in[5].n1 ui_in[5].t0 212.081
R3814 ui_in[5].n6 ui_in[5].t18 212.081
R3815 ui_in[5].n0 ui_in[5].t14 212.081
R3816 ui_in[5].n11 ui_in[5].t16 212.081
R3817 ui_in[5].n17 ui_in[5].t11 212.081
R3818 ui_in[5].n12 ui_in[5].t12 212.081
R3819 ui_in[5].n13 ui_in[5].t15 212.081
R3820 ui_in[5] ui_in[5].n14 163.264
R3821 ui_in[5].n16 ui_in[5].n15 152
R3822 ui_in[5].n19 ui_in[5].n18 152
R3823 ui_in[5].n10 ui_in[5].n9 152
R3824 ui_in[5].n8 ui_in[5].n7 152
R3825 ui_in[5].n5 ui_in[5].n4 152
R3826 ui_in[5] ui_in[5].n3 152
R3827 ui_in[5].n2 ui_in[5].t9 139.78
R3828 ui_in[5].n1 ui_in[5].t10 139.78
R3829 ui_in[5].n6 ui_in[5].t8 139.78
R3830 ui_in[5].n0 ui_in[5].t5 139.78
R3831 ui_in[5].n11 ui_in[5].t7 139.78
R3832 ui_in[5].n17 ui_in[5].t2 139.78
R3833 ui_in[5].n12 ui_in[5].t3 139.78
R3834 ui_in[5].n13 ui_in[5].t6 139.78
R3835 ui_in[5].n24 ui_in[5].t17 120.23
R3836 ui_in[5].n24 ui_in[5].t13 120.228
R3837 ui_in[5].n21 ui_in[5].t4 118.061
R3838 ui_in[5].n21 ui_in[5].t1 118.058
R3839 ui_in[5].n3 ui_in[5].n2 30.6732
R3840 ui_in[5].n3 ui_in[5].n1 30.6732
R3841 ui_in[5].n5 ui_in[5].n1 30.6732
R3842 ui_in[5].n6 ui_in[5].n5 30.6732
R3843 ui_in[5].n7 ui_in[5].n6 30.6732
R3844 ui_in[5].n7 ui_in[5].n0 30.6732
R3845 ui_in[5].n10 ui_in[5].n0 30.6732
R3846 ui_in[5].n11 ui_in[5].n10 30.6732
R3847 ui_in[5].n18 ui_in[5].n11 30.6732
R3848 ui_in[5].n18 ui_in[5].n17 30.6732
R3849 ui_in[5].n17 ui_in[5].n16 30.6732
R3850 ui_in[5].n16 ui_in[5].n12 30.6732
R3851 ui_in[5].n14 ui_in[5].n12 30.6732
R3852 ui_in[5].n14 ui_in[5].n13 30.6732
R3853 ui_in[5].n4 ui_in[5] 21.5045
R3854 ui_in[5].n8 ui_in[5] 19.4565
R3855 ui_in[5].n9 ui_in[5] 17.4085
R3856 ui_in[5].n15 ui_in[5] 13.3125
R3857 ui_in[5].n20 ui_in[5].n19 13.0565
R3858 ui_in[5].n15 ui_in[5] 10.2405
R3859 ui_in[5].n19 ui_in[5] 8.1925
R3860 ui_in[5].n9 ui_in[5] 6.1445
R3861 ui_in[5] ui_in[5].n8 4.0965
R3862 ui_in[5].n23 ui_in[5].n20 3.2054
R3863 ui_in[5].n20 ui_in[5] 2.3045
R3864 ui_in[5].n4 ui_in[5] 2.0485
R3865 ui_in[5].n22 ui_in[5].n21 0.528909
R3866 ui_in[5].n25 ui_in[5].n24 0.506182
R3867 ui_in[5].n26 ui_in[5].n25 0.42675
R3868 ui_in[5].n26 ui_in[5].n23 0.342556
R3869 ui_in[5].n23 ui_in[5].n22 0.3415
R3870 ui_in[5].n25 ui_in[5] 0.170955
R3871 ui_in[5].n22 ui_in[5] 0.148227
R3872 ui_in[5] ui_in[5].n26 0.01225
R3873 ua[0].n4 ua[0].t3 223.565
R3874 ua[0].n7 ua[0].t2 223.565
R3875 ua[0].n0 ua[0].t4 118.769
R3876 ua[0].n3 ua[0].t7 118.621
R3877 ua[0].n2 ua[0].t5 118.005
R3878 ua[0].n1 ua[0].t6 118.005
R3879 ua[0].n0 ua[0].t8 118.005
R3880 ua[0].n6 ua[0].n5 90.2112
R3881 ua[0].n6 ua[0].n4 66.2405
R3882 ua[0].n7 ua[0].n6 63.2157
R3883 ua[0].n5 ua[0].t1 17.4005
R3884 ua[0].n5 ua[0].t0 17.4005
R3885 ua[0].n8 ua[0].n4 5.54823
R3886 ua[0].n8 ua[0].n7 5.18686
R3887 ua[0].n9 ua[0] 4.4438
R3888 ua[0] ua[0].n3 2.77717
R3889 ua[0].n1 ua[0].n0 2.66195
R3890 ua[0].n3 ua[0].n2 1.71868
R3891 ua[0].n2 ua[0].n1 0.764886
R3892 ua[0].n9 ua[0] 0.490406
R3893 ua[0] ua[0].n8 0.244818
R3894 ua[0].n10 ua[0] 0.0992
R3895 ua[0].n10 ua[0] 0.0416941
R3896 ua[0] ua[0].n10 0.0197067
R3897 ua[0] ua[0].n9 0.0129412
R3898 ui_in[1].n2 ui_in[1].t8 212.081
R3899 ui_in[1].n1 ui_in[1].t11 212.081
R3900 ui_in[1].n6 ui_in[1].t7 212.081
R3901 ui_in[1].n0 ui_in[1].t4 212.081
R3902 ui_in[1].n11 ui_in[1].t10 212.081
R3903 ui_in[1].n17 ui_in[1].t6 212.081
R3904 ui_in[1].n12 ui_in[1].t9 212.081
R3905 ui_in[1].n13 ui_in[1].t5 212.081
R3906 ui_in[1] ui_in[1].n14 163.264
R3907 ui_in[1].n16 ui_in[1].n15 152
R3908 ui_in[1].n19 ui_in[1].n18 152
R3909 ui_in[1].n10 ui_in[1].n9 152
R3910 ui_in[1].n8 ui_in[1].n7 152
R3911 ui_in[1].n5 ui_in[1].n4 152
R3912 ui_in[1] ui_in[1].n3 152
R3913 ui_in[1].n2 ui_in[1].t18 139.78
R3914 ui_in[1].n1 ui_in[1].t2 139.78
R3915 ui_in[1].n6 ui_in[1].t17 139.78
R3916 ui_in[1].n0 ui_in[1].t12 139.78
R3917 ui_in[1].n11 ui_in[1].t1 139.78
R3918 ui_in[1].n17 ui_in[1].t16 139.78
R3919 ui_in[1].n12 ui_in[1].t19 139.78
R3920 ui_in[1].n13 ui_in[1].t13 139.78
R3921 ui_in[1].n24 ui_in[1].t0 120.23
R3922 ui_in[1].n24 ui_in[1].t3 120.228
R3923 ui_in[1].n21 ui_in[1].t14 118.061
R3924 ui_in[1].n21 ui_in[1].t15 118.058
R3925 ui_in[1].n3 ui_in[1].n2 30.6732
R3926 ui_in[1].n3 ui_in[1].n1 30.6732
R3927 ui_in[1].n5 ui_in[1].n1 30.6732
R3928 ui_in[1].n6 ui_in[1].n5 30.6732
R3929 ui_in[1].n7 ui_in[1].n6 30.6732
R3930 ui_in[1].n7 ui_in[1].n0 30.6732
R3931 ui_in[1].n10 ui_in[1].n0 30.6732
R3932 ui_in[1].n11 ui_in[1].n10 30.6732
R3933 ui_in[1].n18 ui_in[1].n11 30.6732
R3934 ui_in[1].n18 ui_in[1].n17 30.6732
R3935 ui_in[1].n17 ui_in[1].n16 30.6732
R3936 ui_in[1].n16 ui_in[1].n12 30.6732
R3937 ui_in[1].n14 ui_in[1].n12 30.6732
R3938 ui_in[1].n14 ui_in[1].n13 30.6732
R3939 ui_in[1].n4 ui_in[1] 21.5045
R3940 ui_in[1].n8 ui_in[1] 19.4565
R3941 ui_in[1].n9 ui_in[1] 17.4085
R3942 ui_in[1].n15 ui_in[1] 13.3125
R3943 ui_in[1].n20 ui_in[1].n19 13.0565
R3944 ui_in[1].n15 ui_in[1] 10.2405
R3945 ui_in[1].n19 ui_in[1] 8.1925
R3946 ui_in[1].n9 ui_in[1] 6.1445
R3947 ui_in[1] ui_in[1].n8 4.0965
R3948 ui_in[1].n23 ui_in[1].n20 3.2054
R3949 ui_in[1].n20 ui_in[1] 2.3045
R3950 ui_in[1].n4 ui_in[1] 2.0485
R3951 ui_in[1].n22 ui_in[1].n21 0.528909
R3952 ui_in[1].n25 ui_in[1].n24 0.506182
R3953 ui_in[1].n26 ui_in[1].n25 0.42675
R3954 ui_in[1].n26 ui_in[1].n23 0.342556
R3955 ui_in[1].n23 ui_in[1].n22 0.3415
R3956 ui_in[1].n25 ui_in[1] 0.170955
R3957 ui_in[1].n22 ui_in[1] 0.148227
R3958 ui_in[1] ui_in[1].n26 0.01225
C0 distortionUnit_3.tgate_1.CTRLB distortionUnit_4.IN 1.62697f
C1 ui_in[2] distortionUnit_3.IN 1.74342f
C2 a_20842_23723# distortionUnit_6.IN 0.763261f
C3 distortionUnit_4.myOpamp_0.INn ui_in[3] 0.254411f
C4 distortionUnit_2.myOpamp_0.INn distortionUnit_2.tgate_1.CTRLB 9.98e-19
C5 distortionUnit_5.IN distortionUnit_6.IN 1.38229f
C6 distortionUnit_7.tgate_1.CTRLB VPWR 4.29808f
C7 a_19680_36146# bufferUnit_0.OUT 0.198383f
C8 distortionUnit_6.myOpamp_0.INn distortionUnit_6.IN 0.503808f
C9 ui_in[7] ua[1] 1.87785f
C10 distortionUnit_3.tgate_1.IN distortionUnit_3.IN 0.820736f
C11 VPWR a_7994_36483# 0.156429f
C12 a_20488_30481# distortionUnit_4.tgate_1.IN 2.35765f
C13 distortionUnit_5.IN ui_in[4] 1.59742f
C14 ui_in[1] distortionUnit_2.myOpamp_0.INn 0.254411f
C15 distortionUnit_0.tgate_1.CTRLB distortionUnit_7.IN 1.62697f
C16 distortionUnit_3.myOpamp_0.INn a_6912_30102# 1.1307f
C17 distortionUnit_5.IN distortionUnit_4.tgate_1.CTRLB 1.6595f
C18 distortionUnit_4.IN ui_in[5] 0.291464f
C19 distortionUnit_5.myOpamp_0.INn distortionUnit_5.tgate_1.CTRLB 9.98e-19
C20 VPWR bufferUnit_0.OUT 15.031599f
C21 VPWR a_20584_23723# 4.82533f
C22 ui_in[0] ui_in[4] 0.089269f
C23 ui_in[5] distortionUnit_6.OUT 1.93164f
C24 ui_in[6] distortionUnit_6.IN 0.255482f
C25 a_8014_30557# a_7756_30557# 1.57848f
C26 distortionUnit_0.tgate_1.IN ui_in[6] 0.795971f
C27 distortionUnit_4.tgate_1.IN a_20746_30481# 0.662032f
C28 a_20488_30481# a_19644_30026# 0.27522f
C29 distortionUnit_7.tgate_1.IN distortionUnit_7.IN 0.820736f
C30 a_7032_23398# distortionUnit_5.IN 0.198383f
C31 distortionUnit_6.IN distortionUnit_5.tgate_1.IN 1.38344f
C32 ui_in[4] ui_in[6] 3.36528f
C33 VPWR a_20842_23723# 0.164659f
C34 distortionUnit_5.tgate_1.CTRLB distortionUnit_6.OUT 0.028102f
C35 distortionUnit_4.tgate_1.IN distortionUnit_4.myOpamp_0.INn 1.8069f
C36 a_8134_23853# a_7876_23853# 1.57848f
C37 VPWR bufferUnit_0.tgate_1.CTRLB 4.31158f
C38 distortionUnit_5.IN VPWR 15.008299f
C39 distortionUnit_6.tgate_1.IN distortionUnit_6.OUT 1.38344f
C40 a_21192_16677# distortionUnit_7.IN 0.763261f
C41 VPWR distortionUnit_6.myOpamp_0.INn 1.37899f
C42 VPWR ui_in[0] 5.34653f
C43 a_20746_30481# a_19644_30026# 1.5318f
C44 a_6908_16352# distortionUnit_0.tgate_1.IN 0.001336f
C45 ui_in[4] distortionUnit_5.tgate_1.IN 0.795971f
C46 ui_in[3] ui_in[4] 3.73034f
C47 distortionUnit_5.myOpamp_0.INn a_7876_23853# 0.849481f
C48 distortionUnit_4.tgate_1.CTRLB ui_in[3] 2.30483f
C49 distortionUnit_7.IN distortionUnit_0.tgate_1.IN 1.38344f
C50 distortionUnit_7.myOpamp_0.INn distortionUnit_7.IN 0.503808f
C51 a_6912_30102# distortionUnit_3.tgate_1.IN 0.001336f
C52 a_20524_36601# a_20782_36601# 1.57848f
C53 distortionUnit_4.myOpamp_0.INn a_19644_30026# 1.1307f
C54 a_8014_30557# distortionUnit_3.IN 0.763261f
C55 distortionUnit_6.tgate_1.CTRLB distortionUnit_6.IN 0.258603f
C56 ui_in[2] ui_in[4] 1.79375f
C57 distortionUnit_6.tgate_1.IN ui_in[5] 0.795971f
C58 ui_in[1] ui_in[5] 0.172407f
C59 distortionUnit_3.myOpamp_0.INn VPWR 0.696996f
C60 a_19740_23268# distortionUnit_6.OUT 1.03e-19
C61 distortionUnit_3.tgate_1.CTRLB distortionUnit_3.sky130_fd_sc_hd__tap_2_0.VPB 0.175567f
C62 distortionUnit_4.IN distortionUnit_3.sky130_fd_sc_hd__tap_2_0.VPB 4.57e-19
C63 VPWR ui_in[6] 5.42902f
C64 a_20524_36601# distortionUnit_2.myOpamp_0.INn 0.849481f
C65 ui_in[1] distortionUnit_2.tgate_1.CTRLB 2.30483f
C66 distortionUnit_0.tgate_1.CTRLB distortionUnit_0.sky130_fd_sc_hd__tap_2_0.VPB 0.175567f
C67 a_20584_23723# a_20842_23723# 1.57848f
C68 a_7032_23398# distortionUnit_5.tgate_1.IN 0.001336f
C69 bufferUnit_0.tgate_1.CTRLB bufferUnit_0.OUT 1.62697f
C70 a_20934_16677# distortionUnit_7.tgate_1.IN 2.35765f
C71 distortionUnit_7.tgate_1.IN ua[1] 1.38344f
C72 ua[1] ua[0] 0.45455f
C73 VPWR distortionUnit_5.tgate_1.IN 7.4736f
C74 VPWR ui_in[3] 5.65932f
C75 a_20584_23723# distortionUnit_6.myOpamp_0.INn 0.849481f
C76 ui_in[0] bufferUnit_0.OUT 1.89522f
C77 VPWR distortionUnit_7.sky130_fd_sc_hd__tap_2_0.VPB 0.274328f
C78 distortionUnit_4.IN ui_in[7] 0.253945f
C79 a_20934_16677# a_21192_16677# 1.57848f
C80 a_6908_16352# VPWR 0.100029f
C81 VPWR ui_in[2] 5.62914f
C82 VPWR distortionUnit_7.IN 12.891001f
C83 ui_in[7] distortionUnit_6.OUT 0.317052f
C84 distortionUnit_4.tgate_1.IN distortionUnit_4.tgate_1.CTRLB 1.18066f
C85 VPWR distortionUnit_6.sky130_fd_sc_hd__tap_2_0.VPB 0.274328f
C86 a_20934_16677# distortionUnit_7.myOpamp_0.INn 0.849481f
C87 distortionUnit_6.myOpamp_0.INn a_20842_23723# 1.23683f
C88 bufferUnit_0.OUT ui_in[6] 0.234969f
C89 distortionUnit_7.tgate_1.CTRLB distortionUnit_7.sky130_fd_sc_hd__tap_2_0.VPB 0.175567f
C90 distortionUnit_2.myOpamp_0.INn distortionUnit_3.IN 0.23705f
C91 ua[1] distortionUnit_7.myOpamp_0.INn 0.005273f
C92 distortionUnit_6.tgate_1.IN a_19740_23268# 0.001336f
C93 VPWR distortionUnit_6.tgate_1.CTRLB 4.49268f
C94 ui_in[0] bufferUnit_0.tgate_1.CTRLB 2.30483f
C95 distortionUnit_3.tgate_1.IN VPWR 6.64827f
C96 a_8014_30557# a_6912_30102# 1.5318f
C97 distortionUnit_4.IN a_20488_30481# 3.11184f
C98 distortionUnit_7.tgate_1.CTRLB distortionUnit_7.IN 0.258603f
C99 ui_in[7] ui_in[5] 2.54379f
C100 distortionUnit_0.tgate_1.CTRLB distortionUnit_0.myOpamp_0.INn 9.98e-19
C101 bufferUnit_0.OUT ui_in[3] 0.284299f
C102 distortionUnit_3.myOpamp_0.INn distortionUnit_5.IN 0.190753f
C103 ua[0] bufferUnit_0.tgate_1.IN 1.32325f
C104 distortionUnit_5.sky130_fd_sc_hd__tap_2_0.VPB distortionUnit_6.IN 4.57e-19
C105 distortionUnit_7.tgate_1.IN a_20090_16222# 0.001336f
C106 VPWR distortionUnit_4.tgate_1.IN 6.29098f
C107 a_7752_16807# distortionUnit_0.tgate_1.IN 2.35765f
C108 ui_in[2] bufferUnit_0.OUT 0.262414f
C109 distortionUnit_5.IN ui_in[6] 0.232865f
C110 a_7736_36483# bufferUnit_0.tgate_1.IN 3.21338f
C111 distortionUnit_3.tgate_1.CTRLB distortionUnit_3.IN 0.258603f
C112 distortionUnit_4.IN distortionUnit_3.IN 1.61854f
C113 ui_in[0] ui_in[6] 0.088028f
C114 distortionUnit_4.IN a_20746_30481# 0.763261f
C115 ui_in[7] ui_in[1] 0.18869f
C116 distortionUnit_5.sky130_fd_sc_hd__tap_2_0.VPB ui_in[4] 0.278876f
C117 distortionUnit_5.IN distortionUnit_5.tgate_1.IN 0.820736f
C118 a_21192_16677# a_20090_16222# 1.5318f
C119 distortionUnit_5.IN ui_in[3] 1.92809f
C120 a_20934_16677# VPWR 4.53263f
C121 distortionUnit_4.IN distortionUnit_4.myOpamp_0.INn 0.503808f
C122 ua[1] VPWR 3.53963f
C123 VPWR a_19644_30026# 0.101675f
C124 distortionUnit_0.tgate_1.IN a_8010_16807# 0.662032f
C125 ui_in[0] ui_in[3] 0.089682f
C126 ui_in[2] bufferUnit_0.tgate_1.CTRLB 0.005276f
C127 distortionUnit_7.myOpamp_0.INn a_20090_16222# 1.1307f
C128 distortionUnit_5.IN ui_in[2] 0.044883f
C129 distortionUnit_0.tgate_1.CTRLB distortionUnit_6.OUT 0.258603f
C130 distortionUnit_3.IN ui_in[5] 0.233538f
C131 VPWR distortionUnit_0.sky130_fd_sc_hd__tap_2_0.VPB 0.274328f
C132 distortionUnit_0.tgate_1.IN distortionUnit_0.myOpamp_0.INn 1.8069f
C133 ui_in[0] ui_in[2] 1.02984f
C134 distortionUnit_2.tgate_1.IN a_20782_36601# 0.662032f
C135 a_8014_30557# VPWR 0.161318f
C136 distortionUnit_2.tgate_1.CTRLB distortionUnit_3.IN 1.65953f
C137 ua[1] distortionUnit_7.tgate_1.CTRLB 1.62697f
C138 distortionUnit_4.myOpamp_0.INn ui_in[5] 0.03372f
C139 ui_in[3] ui_in[6] 0.166581f
C140 distortionUnit_5.myOpamp_0.INn distortionUnit_6.IN 0.005273f
C141 VPWR a_7752_16807# 4.63532f
C142 a_6892_36028# distortionUnit_3.IN 3.64e-19
C143 distortionUnit_2.tgate_1.IN distortionUnit_2.myOpamp_0.INn 1.8069f
C144 distortionUnit_2.tgate_1.CTRLB distortionUnit_2.sky130_fd_sc_hd__tap_2_0.VPB 0.175567f
C145 VPWR distortionUnit_5.sky130_fd_sc_hd__tap_2_0.VPB 0.274328f
C146 distortionUnit_6.myOpamp_0.INn distortionUnit_6.tgate_1.CTRLB 9.98e-19
C147 distortionUnit_3.myOpamp_0.INn ui_in[2] 0.254411f
C148 ui_in[2] ui_in[6] 0.085933f
C149 ui_in[1] distortionUnit_3.IN 1.92857f
C150 a_20782_36601# a_19680_36146# 1.5318f
C151 distortionUnit_7.IN ui_in[6] 1.90243f
C152 distortionUnit_5.myOpamp_0.INn ui_in[4] 0.254411f
C153 ui_in[1] distortionUnit_2.sky130_fd_sc_hd__tap_2_0.VPB 0.278876f
C154 distortionUnit_5.IN distortionUnit_4.tgate_1.IN 1.38344f
C155 distortionUnit_3.myOpamp_0.INn distortionUnit_3.tgate_1.IN 1.8069f
C156 VPWR bufferUnit_0.tgate_1.IN 6.64302f
C157 VPWR a_8010_16807# 0.156762f
C158 distortionUnit_2.myOpamp_0.INn a_19680_36146# 1.1307f
C159 distortionUnit_6.IN distortionUnit_6.OUT 1.3678f
C160 ui_in[2] ui_in[3] 3.92737f
C161 a_20090_16222# VPWR 0.100029f
C162 VPWR a_20782_36601# 0.164599f
C163 distortionUnit_0.tgate_1.IN distortionUnit_6.OUT 0.820736f
C164 a_8134_23853# a_7032_23398# 1.5318f
C165 VPWR distortionUnit_0.myOpamp_0.INn 0.877451f
C166 distortionUnit_4.IN ui_in[4] 0.261488f
C167 distortionUnit_4.IN distortionUnit_4.tgate_1.CTRLB 0.258603f
C168 ua[0] a_6892_36028# 0.198383f
C169 a_8134_23853# VPWR 0.193581f
C170 VPWR distortionUnit_2.myOpamp_0.INn 0.866079f
C171 ui_in[4] distortionUnit_6.OUT 0.043613f
C172 distortionUnit_5.IN a_19644_30026# 5.62e-21
C173 distortionUnit_5.myOpamp_0.INn a_7032_23398# 1.1307f
C174 ui_in[5] distortionUnit_6.IN 1.32192f
C175 bufferUnit_0.tgate_1.IN a_7994_36483# 1.89701f
C176 a_7736_36483# a_6892_36028# 0.27522f
C177 distortionUnit_4.tgate_1.CTRLB distortionUnit_4.sky130_fd_sc_hd__tap_2_0.VPB 0.175567f
C178 distortionUnit_5.myOpamp_0.INn VPWR 1.83689f
C179 distortionUnit_3.tgate_1.IN ui_in[2] 0.795971f
C180 bufferUnit_0.tgate_1.IN bufferUnit_0.OUT 1.38344f
C181 ui_in[4] ui_in[5] 3.90346f
C182 distortionUnit_6.tgate_1.CTRLB distortionUnit_6.sky130_fd_sc_hd__tap_2_0.VPB 0.175567f
C183 distortionUnit_4.tgate_1.IN ui_in[3] 0.795971f
C184 distortionUnit_5.tgate_1.CTRLB distortionUnit_6.IN 1.62697f
C185 distortionUnit_2.tgate_1.IN distortionUnit_2.tgate_1.CTRLB 1.18066f
C186 a_20782_36601# bufferUnit_0.OUT 0.763261f
C187 distortionUnit_3.tgate_1.CTRLB VPWR 4.37241f
C188 distortionUnit_4.IN VPWR 15.4213f
C189 ui_in[7] distortionUnit_3.IN 0.240454f
C190 distortionUnit_6.tgate_1.IN distortionUnit_6.IN 0.820736f
C191 a_7756_30557# distortionUnit_3.IN 3.11184f
C192 VPWR distortionUnit_6.OUT 13.9941f
C193 distortionUnit_2.myOpamp_0.INn bufferUnit_0.OUT 0.503808f
C194 distortionUnit_0.sky130_fd_sc_hd__tap_2_0.VPB ui_in[6] 0.278876f
C195 VPWR distortionUnit_4.sky130_fd_sc_hd__tap_2_0.VPB 0.274328f
C196 distortionUnit_3.myOpamp_0.INn a_8014_30557# 1.23683f
C197 distortionUnit_5.tgate_1.CTRLB ui_in[4] 2.30483f
C198 ui_in[1] distortionUnit_2.tgate_1.IN 0.795971f
C199 bufferUnit_0.tgate_1.IN bufferUnit_0.tgate_1.CTRLB 1.18503f
C200 ui_in[1] ui_in[4] 0.174472f
C201 ua[1] distortionUnit_7.sky130_fd_sc_hd__tap_2_0.VPB 4.57e-19
C202 ui_in[0] bufferUnit_0.tgate_1.IN 0.796592f
C203 a_19740_23268# distortionUnit_6.IN 0.198383f
C204 VPWR ui_in[5] 5.68023f
C205 a_20488_30481# a_20746_30481# 1.57848f
C206 a_20934_16677# distortionUnit_7.IN 3.11184f
C207 ua[1] distortionUnit_7.IN 1.3678f
C208 a_8134_23853# distortionUnit_5.IN 0.763261f
C209 VPWR distortionUnit_2.tgate_1.CTRLB 4.40905f
C210 distortionUnit_7.tgate_1.IN ui_in[7] 0.795971f
C211 a_20488_30481# distortionUnit_4.myOpamp_0.INn 0.849481f
C212 VPWR a_6892_36028# 0.102228f
C213 distortionUnit_7.IN distortionUnit_0.sky130_fd_sc_hd__tap_2_0.VPB 4.57e-19
C214 distortionUnit_5.tgate_1.CTRLB VPWR 4.58465f
C215 distortionUnit_5.myOpamp_0.INn distortionUnit_5.IN 0.503808f
C216 distortionUnit_3.IN distortionUnit_2.sky130_fd_sc_hd__tap_2_0.VPB 0.001804f
C217 a_6908_16352# a_7752_16807# 0.27522f
C218 VPWR distortionUnit_6.tgate_1.IN 7.26461f
C219 VPWR ui_in[1] 5.30897f
C220 distortionUnit_0.myOpamp_0.INn ui_in[6] 0.254411f
C221 a_8014_30557# distortionUnit_3.tgate_1.IN 0.662032f
C222 a_6912_30102# a_7756_30557# 0.27522f
C223 ui_in[7] distortionUnit_6.IN 0.267407f
C224 distortionUnit_4.myOpamp_0.INn a_20746_30481# 1.23683f
C225 bufferUnit_0.OUT ui_in[5] 0.238698f
C226 distortionUnit_3.tgate_1.CTRLB distortionUnit_5.IN 0.028918f
C227 distortionUnit_4.IN distortionUnit_5.IN 1.3678f
C228 ui_in[7] distortionUnit_7.myOpamp_0.INn 0.254411f
C229 distortionUnit_3.IN bufferUnit_0.sky130_fd_sc_hd__tap_2_0.VPB 0.001611f
C230 distortionUnit_4.tgate_1.IN a_19644_30026# 0.001336f
C231 a_7994_36483# a_6892_36028# 1.5318f
C232 distortionUnit_2.tgate_1.CTRLB bufferUnit_0.OUT 0.258603f
C233 a_6908_16352# a_8010_16807# 1.5318f
C234 VPWR a_19740_23268# 0.120584f
C235 distortionUnit_5.IN distortionUnit_4.sky130_fd_sc_hd__tap_2_0.VPB 0.001804f
C236 a_20524_36601# distortionUnit_2.tgate_1.IN 2.35765f
C237 ui_in[7] ui_in[4] 0.089626f
C238 distortionUnit_6.myOpamp_0.INn distortionUnit_6.OUT 0.260919f
C239 a_8134_23853# distortionUnit_5.tgate_1.IN 0.662032f
C240 a_7032_23398# a_7876_23853# 0.27522f
C241 distortionUnit_2.myOpamp_0.INn ui_in[3] 0.058805f
C242 a_20090_16222# distortionUnit_7.IN 0.198383f
C243 a_6908_16352# distortionUnit_0.myOpamp_0.INn 1.1307f
C244 VPWR a_7876_23853# 5.38803f
C245 VPWR distortionUnit_3.sky130_fd_sc_hd__tap_2_0.VPB 0.274328f
C246 distortionUnit_3.myOpamp_0.INn distortionUnit_3.tgate_1.CTRLB 9.98e-19
C247 distortionUnit_3.myOpamp_0.INn distortionUnit_4.IN 0.005273f
C248 a_20584_23723# distortionUnit_6.tgate_1.IN 2.35765f
C249 distortionUnit_5.myOpamp_0.INn distortionUnit_5.tgate_1.IN 1.8069f
C250 ui_in[1] bufferUnit_0.OUT 1.59433f
C251 distortionUnit_7.IN distortionUnit_0.myOpamp_0.INn 0.005273f
C252 distortionUnit_5.IN ui_in[5] 0.337455f
C253 distortionUnit_4.IN ui_in[6] 0.244964f
C254 distortionUnit_6.myOpamp_0.INn ui_in[5] 0.254411f
C255 ui_in[0] ui_in[5] 0.087906f
C256 a_20524_36601# a_19680_36146# 0.27522f
C257 ui_in[6] distortionUnit_6.OUT 1.58548f
C258 a_6912_30102# distortionUnit_3.IN 0.198383f
C259 distortionUnit_4.IN ui_in[3] 1.31839f
C260 distortionUnit_5.tgate_1.CTRLB distortionUnit_5.IN 0.258603f
C261 ui_in[7] VPWR 5.46148f
C262 a_20584_23723# a_19740_23268# 0.27522f
C263 distortionUnit_6.tgate_1.IN a_20842_23723# 0.662032f
C264 a_7756_30557# VPWR 4.6075f
C265 distortionUnit_2.tgate_1.IN distortionUnit_3.IN 1.38344f
C266 VPWR a_20524_36601# 4.64125f
C267 distortionUnit_4.sky130_fd_sc_hd__tap_2_0.VPB ui_in[3] 0.278876f
C268 distortionUnit_3.IN ui_in[4] 0.234366f
C269 ui_in[5] ui_in[6] 3.7149f
C270 distortionUnit_3.tgate_1.CTRLB ui_in[2] 2.30483f
C271 distortionUnit_4.IN ui_in[2] 1.89891f
C272 distortionUnit_6.tgate_1.IN distortionUnit_6.myOpamp_0.INn 1.8069f
C273 ui_in[0] ui_in[1] 4.72532f
C274 distortionUnit_0.tgate_1.CTRLB distortionUnit_0.tgate_1.IN 1.18066f
C275 a_6908_16352# distortionUnit_6.OUT 0.198383f
C276 ua[0] a_7736_36483# 3.11184f
C277 ui_in[7] distortionUnit_7.tgate_1.CTRLB 2.30483f
C278 distortionUnit_7.IN distortionUnit_6.OUT 1.3678f
C279 a_20842_23723# a_19740_23268# 1.5318f
C280 a_20934_16677# a_20090_16222# 0.27522f
C281 distortionUnit_7.tgate_1.IN a_21192_16677# 0.662032f
C282 VPWR a_20488_30481# 4.57345f
C283 distortionUnit_3.tgate_1.CTRLB distortionUnit_3.tgate_1.IN 1.18066f
C284 ui_in[3] ui_in[5] 2.18372f
C285 distortionUnit_4.IN distortionUnit_3.tgate_1.IN 1.38344f
C286 a_19680_36146# distortionUnit_3.IN 5.62e-21
C287 distortionUnit_4.myOpamp_0.INn distortionUnit_4.tgate_1.CTRLB 9.98e-19
C288 distortionUnit_6.sky130_fd_sc_hd__tap_2_0.VPB distortionUnit_6.OUT 0.001873f
C289 distortionUnit_6.tgate_1.CTRLB distortionUnit_6.OUT 1.66142f
C290 distortionUnit_6.myOpamp_0.INn a_19740_23268# 1.1307f
C291 distortionUnit_7.tgate_1.IN distortionUnit_7.myOpamp_0.INn 1.8069f
C292 ui_in[2] ui_in[5] 0.086037f
C293 ui_in[1] ui_in[6] 0.17014f
C294 ui_in[7] bufferUnit_0.OUT 0.24347f
C295 distortionUnit_5.IN a_7876_23853# 3.11184f
C296 distortionUnit_5.IN distortionUnit_3.sky130_fd_sc_hd__tap_2_0.VPB 0.001206f
C297 a_20524_36601# bufferUnit_0.OUT 3.11184f
C298 distortionUnit_5.tgate_1.CTRLB distortionUnit_5.tgate_1.IN 1.18066f
C299 VPWR distortionUnit_3.IN 14.9278f
C300 distortionUnit_6.sky130_fd_sc_hd__tap_2_0.VPB ui_in[5] 0.278876f
C301 VPWR a_20746_30481# 0.156113f
C302 a_7752_16807# a_8010_16807# 1.57848f
C303 distortionUnit_4.IN distortionUnit_4.tgate_1.IN 0.820736f
C304 distortionUnit_6.tgate_1.CTRLB ui_in[5] 2.30483f
C305 VPWR distortionUnit_2.sky130_fd_sc_hd__tap_2_0.VPB 0.274328f
C306 ui_in[1] ui_in[3] 1.03886f
C307 distortionUnit_7.myOpamp_0.INn a_21192_16677# 1.23683f
C308 VPWR distortionUnit_4.myOpamp_0.INn 0.577656f
C309 a_7752_16807# distortionUnit_0.myOpamp_0.INn 0.849481f
C310 distortionUnit_0.tgate_1.CTRLB VPWR 4.4067f
C311 ui_in[1] ui_in[2] 4.51989f
C312 distortionUnit_5.IN ui_in[7] 0.238801f
C313 VPWR bufferUnit_0.sky130_fd_sc_hd__tap_2_0.VPB 0.274803f
C314 ui_in[4] distortionUnit_6.IN 1.90075f
C315 distortionUnit_4.IN a_19644_30026# 0.198383f
C316 ui_in[7] distortionUnit_6.myOpamp_0.INn 0.030058f
C317 ui_in[7] ui_in[0] 0.089842f
C318 distortionUnit_6.tgate_1.IN distortionUnit_6.tgate_1.CTRLB 1.18066f
C319 distortionUnit_7.tgate_1.IN VPWR 6.25246f
C320 bufferUnit_0.OUT distortionUnit_3.IN 1.3678f
C321 distortionUnit_0.myOpamp_0.INn a_8010_16807# 1.23683f
C322 VPWR ua[0] 20.5546f
C323 a_7876_23853# distortionUnit_5.tgate_1.IN 2.35765f
C324 distortionUnit_3.myOpamp_0.INn a_7756_30557# 0.849481f
C325 VPWR a_7736_36483# 4.57503f
C326 distortionUnit_2.myOpamp_0.INn a_20782_36601# 1.23683f
C327 ui_in[7] ui_in[6] 7.30655f
C328 ui_in[2] distortionUnit_3.sky130_fd_sc_hd__tap_2_0.VPB 0.278876f
C329 a_21192_16677# VPWR 0.148886f
C330 distortionUnit_2.tgate_1.IN a_19680_36146# 0.001336f
C331 distortionUnit_7.tgate_1.IN distortionUnit_7.tgate_1.CTRLB 1.18066f
C332 a_7752_16807# distortionUnit_6.OUT 3.11184f
C333 a_6912_30102# VPWR 0.124672f
C334 distortionUnit_5.sky130_fd_sc_hd__tap_2_0.VPB distortionUnit_6.OUT 0.001173f
C335 bufferUnit_0.OUT bufferUnit_0.sky130_fd_sc_hd__tap_2_0.VPB 4.57e-19
C336 VPWR distortionUnit_6.IN 14.791201f
C337 VPWR distortionUnit_0.tgate_1.IN 6.91249f
C338 bufferUnit_0.tgate_1.CTRLB distortionUnit_3.IN 0.040054f
C339 distortionUnit_5.IN distortionUnit_3.IN 0.185605f
C340 ua[0] a_7994_36483# 0.763261f
C341 distortionUnit_7.myOpamp_0.INn VPWR 0.533126f
C342 ui_in[7] ui_in[3] 0.184684f
C343 distortionUnit_5.myOpamp_0.INn a_8134_23853# 1.23683f
C344 ui_in[7] distortionUnit_7.sky130_fd_sc_hd__tap_2_0.VPB 0.278876f
C345 VPWR distortionUnit_2.tgate_1.IN 6.88903f
C346 ui_in[0] distortionUnit_3.IN 0.062373f
C347 a_7736_36483# a_7994_36483# 1.57848f
C348 ua[0] bufferUnit_0.OUT 1.3678f
C349 VPWR ui_in[4] 5.66885f
C350 ui_in[7] ui_in[2] 0.086999f
C351 VPWR distortionUnit_4.tgate_1.CTRLB 4.30804f
C352 distortionUnit_5.IN distortionUnit_4.myOpamp_0.INn 0.236699f
C353 a_8010_16807# distortionUnit_6.OUT 0.763261f
C354 ui_in[7] distortionUnit_7.IN 1.33097f
C355 distortionUnit_7.myOpamp_0.INn distortionUnit_7.tgate_1.CTRLB 9.98e-19
C356 bufferUnit_0.tgate_1.CTRLB bufferUnit_0.sky130_fd_sc_hd__tap_2_0.VPB 0.175567f
C357 distortionUnit_3.myOpamp_0.INn distortionUnit_3.IN 0.503808f
C358 distortionUnit_0.myOpamp_0.INn distortionUnit_6.OUT 0.503808f
C359 VPWR a_19680_36146# 0.138823f
C360 distortionUnit_3.IN ui_in[6] 0.234443f
C361 ui_in[0] bufferUnit_0.sky130_fd_sc_hd__tap_2_0.VPB 0.278876f
C362 a_7756_30557# distortionUnit_3.tgate_1.IN 2.35765f
C363 distortionUnit_5.tgate_1.CTRLB distortionUnit_5.sky130_fd_sc_hd__tap_2_0.VPB 0.175567f
C364 a_20584_23723# distortionUnit_6.IN 3.11184f
C365 ua[0] bufferUnit_0.tgate_1.CTRLB 0.258603f
C366 a_7032_23398# VPWR 0.185809f
C367 distortionUnit_5.myOpamp_0.INn distortionUnit_6.OUT 0.182465f
C368 distortionUnit_2.tgate_1.IN bufferUnit_0.OUT 0.820736f
C369 distortionUnit_3.IN ui_in[3] 1.11357f
C370 ui_in[0] ua[0] 1.3091f
C371 bufferUnit_0.tgate_1.IN a_6892_36028# 1.13204f
C372 distortionUnit_0.tgate_1.CTRLB ui_in[6] 2.30483f
C373 bufferUnit_0.OUT ui_in[4] 0.236467f
C374 ua[1] VGND 20.273489f
C375 ui_in[7] VGND 30.44768f
C376 ui_in[6] VGND 28.305063f
C377 ui_in[5] VGND 28.04585f
C378 ui_in[4] VGND 24.38101f
C379 ui_in[3] VGND 24.551018f
C380 ui_in[2] VGND 21.405066f
C381 ui_in[1] VGND 21.530848f
C382 ua[0] VGND 60.802273f
C383 ui_in[0] VGND 20.53937f
C384 VPWR VGND -0.245118p
C385 distortionUnit_7.tgate_1.CTRLB VGND 4.90752f
C386 a_20090_16222# VGND 5.77906f
C387 a_21192_16677# VGND 1.79918f
C388 distortionUnit_7.myOpamp_0.INn VGND 8.745749f
C389 distortionUnit_7.tgate_1.IN VGND 2.7889f
C390 a_20934_16677# VGND 4.02935f
C391 distortionUnit_0.tgate_1.CTRLB VGND 4.9219f
C392 a_6908_16352# VGND 5.75903f
C393 a_8010_16807# VGND 1.78029f
C394 distortionUnit_0.myOpamp_0.INn VGND 8.475241f
C395 distortionUnit_0.tgate_1.IN VGND 2.55922f
C396 a_7752_16807# VGND 3.58914f
C397 distortionUnit_7.IN VGND 14.596201f
C398 distortionUnit_6.tgate_1.CTRLB VGND 4.86653f
C399 a_19740_23268# VGND 5.71244f
C400 a_20842_23723# VGND 1.74561f
C401 distortionUnit_6.myOpamp_0.INn VGND 8.006411f
C402 distortionUnit_6.tgate_1.IN VGND 2.46277f
C403 a_20584_23723# VGND 3.11162f
C404 distortionUnit_5.tgate_1.CTRLB VGND 4.79417f
C405 a_7032_23398# VGND 5.62744f
C406 a_8134_23853# VGND 1.69448f
C407 distortionUnit_5.myOpamp_0.INn VGND 8.00655f
C408 distortionUnit_5.tgate_1.IN VGND 2.42202f
C409 a_7876_23853# VGND 2.82463f
C410 distortionUnit_6.OUT VGND 30.3326f
C411 distortionUnit_6.IN VGND 13.4661f
C412 distortionUnit_4.tgate_1.CTRLB VGND 4.89068f
C413 a_19644_30026# VGND 5.73711f
C414 a_20746_30481# VGND 1.75741f
C415 distortionUnit_4.myOpamp_0.INn VGND 8.0762f
C416 distortionUnit_4.tgate_1.IN VGND 2.55307f
C417 a_20488_30481# VGND 3.28069f
C418 distortionUnit_3.tgate_1.CTRLB VGND 4.85582f
C419 a_6912_30102# VGND 5.69131f
C420 a_8014_30557# VGND 1.73604f
C421 distortionUnit_3.myOpamp_0.INn VGND 8.0678f
C422 distortionUnit_3.tgate_1.IN VGND 2.49844f
C423 a_7756_30557# VGND 3.01493f
C424 distortionUnit_5.IN VGND 37.727688f
C425 distortionUnit_4.IN VGND 13.2873f
C426 distortionUnit_2.tgate_1.CTRLB VGND 4.82872f
C427 a_19680_36146# VGND 5.66154f
C428 a_20782_36601# VGND 1.72068f
C429 distortionUnit_2.myOpamp_0.INn VGND 7.96703f
C430 distortionUnit_2.tgate_1.IN VGND 2.47812f
C431 a_20524_36601# VGND 2.92111f
C432 bufferUnit_0.tgate_1.CTRLB VGND 4.88605f
C433 a_6892_36028# VGND 5.73517f
C434 a_7994_36483# VGND 1.75688f
C435 bufferUnit_0.tgate_1.IN VGND 5.32069f
C436 a_7736_36483# VGND 3.2716f
C437 distortionUnit_3.IN VGND 29.748499f
C438 bufferUnit_0.OUT VGND 13.1831f
C439 distortionUnit_7.sky130_fd_sc_hd__tap_2_0.VPB VGND 1.14309f
C440 distortionUnit_0.sky130_fd_sc_hd__tap_2_0.VPB VGND 1.14329f
C441 distortionUnit_6.sky130_fd_sc_hd__tap_2_0.VPB VGND 1.14329f
C442 distortionUnit_5.sky130_fd_sc_hd__tap_2_0.VPB VGND 1.14329f
C443 distortionUnit_4.sky130_fd_sc_hd__tap_2_0.VPB VGND 1.14329f
C444 distortionUnit_3.sky130_fd_sc_hd__tap_2_0.VPB VGND 1.14329f
C445 distortionUnit_2.sky130_fd_sc_hd__tap_2_0.VPB VGND 1.14329f
C446 bufferUnit_0.sky130_fd_sc_hd__tap_2_0.VPB VGND 1.14329f
C447 ui_in[1].t10 VGND 0.012664f
C448 ui_in[1].t1 VGND 0.007463f
C449 ui_in[1].t4 VGND 0.012664f
C450 ui_in[1].t12 VGND 0.007463f
C451 ui_in[1].n0 VGND 0.018264f
C452 ui_in[1].t7 VGND 0.012664f
C453 ui_in[1].t17 VGND 0.007463f
C454 ui_in[1].t11 VGND 0.012664f
C455 ui_in[1].t2 VGND 0.007463f
C456 ui_in[1].n1 VGND 0.018264f
C457 ui_in[1].t8 VGND 0.012664f
C458 ui_in[1].t18 VGND 0.007463f
C459 ui_in[1].n2 VGND 0.01707f
C460 ui_in[1].n3 VGND 0.008358f
C461 ui_in[1].n4 VGND 0.006935f
C462 ui_in[1].n5 VGND 0.008358f
C463 ui_in[1].n6 VGND 0.018264f
C464 ui_in[1].n7 VGND 0.008358f
C465 ui_in[1].n8 VGND 0.006935f
C466 ui_in[1].n9 VGND 0.006935f
C467 ui_in[1].n10 VGND 0.008358f
C468 ui_in[1].n11 VGND 0.018264f
C469 ui_in[1].t6 VGND 0.012664f
C470 ui_in[1].t16 VGND 0.007463f
C471 ui_in[1].t9 VGND 0.012664f
C472 ui_in[1].t19 VGND 0.007463f
C473 ui_in[1].n12 VGND 0.018264f
C474 ui_in[1].t5 VGND 0.012664f
C475 ui_in[1].t13 VGND 0.007463f
C476 ui_in[1].n13 VGND 0.01707f
C477 ui_in[1].n14 VGND 0.00893f
C478 ui_in[1].n15 VGND 0.006935f
C479 ui_in[1].n16 VGND 0.008358f
C480 ui_in[1].n17 VGND 0.018264f
C481 ui_in[1].n18 VGND 0.008358f
C482 ui_in[1].n19 VGND 0.006257f
C483 ui_in[1].n20 VGND 0.42528f
C484 ui_in[1].t14 VGND 0.137801f
C485 ui_in[1].t15 VGND 0.137799f
C486 ui_in[1].n21 VGND 0.797557f
C487 ui_in[1].n22 VGND 0.523381f
C488 ui_in[1].n23 VGND 2.78149f
C489 ui_in[1].t0 VGND 0.141499f
C490 ui_in[1].t3 VGND 0.141497f
C491 ui_in[1].n24 VGND 0.780809f
C492 ui_in[1].n25 VGND 0.529164f
C493 ui_in[1].n26 VGND 1.47086f
C494 ua[0].t4 VGND 0.044976f
C495 ua[0].t8 VGND 0.044828f
C496 ua[0].n0 VGND 0.055526f
C497 ua[0].t6 VGND 0.044828f
C498 ua[0].n1 VGND 0.032759f
C499 ua[0].t5 VGND 0.044828f
C500 ua[0].n2 VGND 0.028433f
C501 ua[0].t7 VGND 0.044943f
C502 ua[0].n3 VGND 0.077958f
C503 ua[0].t3 VGND 0.010295f
C504 ua[0].n4 VGND 0.039777f
C505 ua[0].t1 VGND 0.002846f
C506 ua[0].t0 VGND 0.002846f
C507 ua[0].n5 VGND 0.009237f
C508 ua[0].n6 VGND 0.056327f
C509 ua[0].t2 VGND 0.010295f
C510 ua[0].n7 VGND 0.029716f
C511 ua[0].n8 VGND 0.3405f
C512 ua[0].n9 VGND 1.30885f
C513 ua[0].n10 VGND 0.274984f
C514 ui_in[5].t16 VGND 0.012772f
C515 ui_in[5].t7 VGND 0.007526f
C516 ui_in[5].t14 VGND 0.012772f
C517 ui_in[5].t5 VGND 0.007526f
C518 ui_in[5].n0 VGND 0.018418f
C519 ui_in[5].t18 VGND 0.012772f
C520 ui_in[5].t8 VGND 0.007526f
C521 ui_in[5].t0 VGND 0.012772f
C522 ui_in[5].t10 VGND 0.007526f
C523 ui_in[5].n1 VGND 0.018418f
C524 ui_in[5].t19 VGND 0.012772f
C525 ui_in[5].t9 VGND 0.007526f
C526 ui_in[5].n2 VGND 0.017214f
C527 ui_in[5].n3 VGND 0.008429f
C528 ui_in[5].n4 VGND 0.006994f
C529 ui_in[5].n5 VGND 0.008429f
C530 ui_in[5].n6 VGND 0.018418f
C531 ui_in[5].n7 VGND 0.008429f
C532 ui_in[5].n8 VGND 0.006994f
C533 ui_in[5].n9 VGND 0.006994f
C534 ui_in[5].n10 VGND 0.008429f
C535 ui_in[5].n11 VGND 0.018418f
C536 ui_in[5].t11 VGND 0.012772f
C537 ui_in[5].t2 VGND 0.007526f
C538 ui_in[5].t12 VGND 0.012772f
C539 ui_in[5].t3 VGND 0.007526f
C540 ui_in[5].n12 VGND 0.018418f
C541 ui_in[5].t15 VGND 0.012772f
C542 ui_in[5].t6 VGND 0.007526f
C543 ui_in[5].n13 VGND 0.017214f
C544 ui_in[5].n14 VGND 0.009006f
C545 ui_in[5].n15 VGND 0.006994f
C546 ui_in[5].n16 VGND 0.008429f
C547 ui_in[5].n17 VGND 0.018418f
C548 ui_in[5].n18 VGND 0.008429f
C549 ui_in[5].n19 VGND 0.00631f
C550 ui_in[5].n20 VGND 0.428882f
C551 ui_in[5].t4 VGND 0.138968f
C552 ui_in[5].t1 VGND 0.138967f
C553 ui_in[5].n21 VGND 0.804313f
C554 ui_in[5].n22 VGND 0.527814f
C555 ui_in[5].n23 VGND 2.80505f
C556 ui_in[5].t17 VGND 0.142697f
C557 ui_in[5].t13 VGND 0.142695f
C558 ui_in[5].n24 VGND 0.787423f
C559 ui_in[5].n25 VGND 0.533646f
C560 ui_in[5].n26 VGND 1.48332f
C561 ui_in[2].t9 VGND 0.011838f
C562 ui_in[2].t15 VGND 0.006976f
C563 ui_in[2].t4 VGND 0.011838f
C564 ui_in[2].t12 VGND 0.006976f
C565 ui_in[2].n0 VGND 0.017073f
C566 ui_in[2].t10 VGND 0.011838f
C567 ui_in[2].t16 VGND 0.006976f
C568 ui_in[2].t1 VGND 0.011838f
C569 ui_in[2].t7 VGND 0.006976f
C570 ui_in[2].n1 VGND 0.017073f
C571 ui_in[2].t5 VGND 0.011838f
C572 ui_in[2].t13 VGND 0.006976f
C573 ui_in[2].n2 VGND 0.015957f
C574 ui_in[2].n3 VGND 0.007813f
C575 ui_in[2].n4 VGND 0.006483f
C576 ui_in[2].n5 VGND 0.007813f
C577 ui_in[2].n6 VGND 0.017073f
C578 ui_in[2].n7 VGND 0.007813f
C579 ui_in[2].n8 VGND 0.006483f
C580 ui_in[2].n9 VGND 0.006483f
C581 ui_in[2].n10 VGND 0.007813f
C582 ui_in[2].n11 VGND 0.017073f
C583 ui_in[2].t3 VGND 0.011838f
C584 ui_in[2].t11 VGND 0.006976f
C585 ui_in[2].t0 VGND 0.011838f
C586 ui_in[2].t6 VGND 0.006976f
C587 ui_in[2].n12 VGND 0.017073f
C588 ui_in[2].t2 VGND 0.011838f
C589 ui_in[2].t8 VGND 0.006976f
C590 ui_in[2].n13 VGND 0.015957f
C591 ui_in[2].n14 VGND 0.008348f
C592 ui_in[2].n15 VGND 0.006483f
C593 ui_in[2].n16 VGND 0.007813f
C594 ui_in[2].n17 VGND 0.017073f
C595 ui_in[2].n18 VGND 0.007813f
C596 ui_in[2].n19 VGND 0.005849f
C597 ui_in[2].n20 VGND 0.39755f
C598 ui_in[2].t18 VGND 0.128816f
C599 ui_in[2].t19 VGND 0.128814f
C600 ui_in[2].n21 VGND 0.745554f
C601 ui_in[2].n22 VGND 0.489254f
C602 ui_in[2].n23 VGND 2.60012f
C603 ui_in[2].t14 VGND 0.132272f
C604 ui_in[2].t17 VGND 0.132271f
C605 ui_in[2].n24 VGND 0.729898f
C606 ui_in[2].n25 VGND 0.494661f
C607 ui_in[2].n26 VGND 1.37496f
C608 ui_in[0].t0 VGND 0.009748f
C609 ui_in[0].t10 VGND 0.005744f
C610 ui_in[0].t17 VGND 0.009748f
C611 ui_in[0].t8 VGND 0.005744f
C612 ui_in[0].n0 VGND 0.014058f
C613 ui_in[0].t14 VGND 0.009748f
C614 ui_in[0].t5 VGND 0.005744f
C615 ui_in[0].t12 VGND 0.009748f
C616 ui_in[0].t3 VGND 0.005744f
C617 ui_in[0].n1 VGND 0.014058f
C618 ui_in[0].t18 VGND 0.009748f
C619 ui_in[0].t9 VGND 0.005744f
C620 ui_in[0].n2 VGND 0.013139f
C621 ui_in[0].n3 VGND 0.006434f
C622 ui_in[0].n4 VGND 0.005338f
C623 ui_in[0].n5 VGND 0.006434f
C624 ui_in[0].n6 VGND 0.014058f
C625 ui_in[0].n7 VGND 0.006434f
C626 ui_in[0].n8 VGND 0.005338f
C627 ui_in[0].n9 VGND 0.005338f
C628 ui_in[0].n10 VGND 0.006434f
C629 ui_in[0].n11 VGND 0.014058f
C630 ui_in[0].t16 VGND 0.009748f
C631 ui_in[0].t7 VGND 0.005744f
C632 ui_in[0].t11 VGND 0.009748f
C633 ui_in[0].t1 VGND 0.005744f
C634 ui_in[0].n12 VGND 0.014058f
C635 ui_in[0].t13 VGND 0.009748f
C636 ui_in[0].t4 VGND 0.005744f
C637 ui_in[0].n13 VGND 0.013139f
C638 ui_in[0].n14 VGND 0.006874f
C639 ui_in[0].n15 VGND 0.005338f
C640 ui_in[0].n16 VGND 0.006434f
C641 ui_in[0].n17 VGND 0.014058f
C642 ui_in[0].n18 VGND 0.006434f
C643 ui_in[0].n19 VGND 0.004816f
C644 ui_in[0].n20 VGND 0.327354f
C645 ui_in[0].t2 VGND 0.106071f
C646 ui_in[0].t6 VGND 0.106069f
C647 ui_in[0].n21 VGND 0.613909f
C648 ui_in[0].n22 VGND 0.402866f
C649 ui_in[0].n23 VGND 2.14101f
C650 ui_in[0].t15 VGND 0.108917f
C651 ui_in[0].t19 VGND 0.108915f
C652 ui_in[0].n24 VGND 0.601018f
C653 ui_in[0].n25 VGND 0.407317f
C654 ui_in[0].n26 VGND 1.13218f
C655 ua[1].n0 VGND 0.043178f
C656 ua[1].t5 VGND 0.001064f
C657 ua[1].t4 VGND 0.001064f
C658 ua[1].n1 VGND 0.002204f
C659 ua[1].t0 VGND 0.003846f
C660 ua[1].n2 VGND 0.030935f
C661 ua[1].n3 VGND 0.028972f
C662 ua[1].t1 VGND 0.003805f
C663 ua[1].n4 VGND 0.030242f
C664 ua[1].n5 VGND 0.097005f
C665 ua[1].n6 VGND 0.043178f
C666 ua[1].t2 VGND 0.001064f
C667 ua[1].t3 VGND 0.001064f
C668 ua[1].n7 VGND 0.002204f
C669 ua[1].t6 VGND 0.003846f
C670 ua[1].n8 VGND 0.030935f
C671 ua[1].n9 VGND 0.028972f
C672 ua[1].t7 VGND 0.003805f
C673 ua[1].n10 VGND 0.030242f
C674 ua[1].n11 VGND 0.075781f
C675 ua[1].n12 VGND 0.199199f
C676 ua[1].n13 VGND 1.7979f
C677 ui_in[7].t8 VGND 0.010065f
C678 ui_in[7].t17 VGND 0.005931f
C679 ui_in[7].t4 VGND 0.010065f
C680 ui_in[7].t14 VGND 0.005931f
C681 ui_in[7].n0 VGND 0.014515f
C682 ui_in[7].t3 VGND 0.010065f
C683 ui_in[7].t13 VGND 0.005931f
C684 ui_in[7].t9 VGND 0.010065f
C685 ui_in[7].t18 VGND 0.005931f
C686 ui_in[7].n1 VGND 0.014515f
C687 ui_in[7].t5 VGND 0.010065f
C688 ui_in[7].t15 VGND 0.005931f
C689 ui_in[7].n2 VGND 0.013566f
C690 ui_in[7].n3 VGND 0.006643f
C691 ui_in[7].n4 VGND 0.005512f
C692 ui_in[7].n5 VGND 0.006643f
C693 ui_in[7].n6 VGND 0.014515f
C694 ui_in[7].n7 VGND 0.006643f
C695 ui_in[7].n8 VGND 0.005512f
C696 ui_in[7].n9 VGND 0.005512f
C697 ui_in[7].n10 VGND 0.006643f
C698 ui_in[7].n11 VGND 0.014515f
C699 ui_in[7].t2 VGND 0.010065f
C700 ui_in[7].t12 VGND 0.005931f
C701 ui_in[7].t6 VGND 0.010065f
C702 ui_in[7].t16 VGND 0.005931f
C703 ui_in[7].n12 VGND 0.014515f
C704 ui_in[7].t1 VGND 0.010065f
C705 ui_in[7].t11 VGND 0.005931f
C706 ui_in[7].n13 VGND 0.013566f
C707 ui_in[7].n14 VGND 0.007098f
C708 ui_in[7].n15 VGND 0.005512f
C709 ui_in[7].n16 VGND 0.006643f
C710 ui_in[7].n17 VGND 0.014515f
C711 ui_in[7].n18 VGND 0.006643f
C712 ui_in[7].n19 VGND 0.004973f
C713 ui_in[7].n20 VGND 0.337994f
C714 ui_in[7].t7 VGND 0.109518f
C715 ui_in[7].t10 VGND 0.109517f
C716 ui_in[7].n21 VGND 0.633864f
C717 ui_in[7].n22 VGND 0.41596f
C718 ui_in[7].n23 VGND 2.2106f
C719 ui_in[7].t19 VGND 0.112457f
C720 ui_in[7].t0 VGND 0.112455f
C721 ui_in[7].n24 VGND 0.620553f
C722 ui_in[7].n25 VGND 0.420556f
C723 ui_in[7].n26 VGND 1.16898f
C724 distortionUnit_5.IN.t0 VGND 0.011149f
C725 distortionUnit_5.IN.n0 VGND 0.04308f
C726 distortionUnit_5.IN.t2 VGND 0.003083f
C727 distortionUnit_5.IN.t3 VGND 0.003083f
C728 distortionUnit_5.IN.n1 VGND 0.010004f
C729 distortionUnit_5.IN.n2 VGND 0.061004f
C730 distortionUnit_5.IN.t1 VGND 0.011149f
C731 distortionUnit_5.IN.n3 VGND 0.032184f
C732 distortionUnit_5.IN.n4 VGND 0.368775f
C733 distortionUnit_5.IN.n5 VGND 0.125118f
C734 distortionUnit_5.IN.t11 VGND 0.003083f
C735 distortionUnit_5.IN.t10 VGND 0.003083f
C736 distortionUnit_5.IN.n6 VGND 0.006386f
C737 distortionUnit_5.IN.t7 VGND 0.011144f
C738 distortionUnit_5.IN.n7 VGND 0.089641f
C739 distortionUnit_5.IN.n8 VGND 0.083951f
C740 distortionUnit_5.IN.t6 VGND 0.011026f
C741 distortionUnit_5.IN.n9 VGND 0.087633f
C742 distortionUnit_5.IN.n10 VGND 0.281094f
C743 distortionUnit_5.IN.n11 VGND 0.125118f
C744 distortionUnit_5.IN.t5 VGND 0.003083f
C745 distortionUnit_5.IN.t4 VGND 0.003083f
C746 distortionUnit_5.IN.n12 VGND 0.006386f
C747 distortionUnit_5.IN.t8 VGND 0.011144f
C748 distortionUnit_5.IN.n13 VGND 0.089641f
C749 distortionUnit_5.IN.n14 VGND 0.083951f
C750 distortionUnit_5.IN.t9 VGND 0.011026f
C751 distortionUnit_5.IN.n15 VGND 0.087633f
C752 distortionUnit_5.IN.n16 VGND 0.219593f
C753 distortionUnit_5.IN.n17 VGND 0.577223f
C754 distortionUnit_5.IN.n18 VGND 5.86744f
C755 distortionUnit_5.IN.t14 VGND 0.04871f
C756 distortionUnit_5.IN.t13 VGND 0.048551f
C757 distortionUnit_5.IN.n19 VGND 0.060137f
C758 distortionUnit_5.IN.t15 VGND 0.048551f
C759 distortionUnit_5.IN.n20 VGND 0.03548f
C760 distortionUnit_5.IN.t16 VGND 0.048551f
C761 distortionUnit_5.IN.n21 VGND 0.030794f
C762 distortionUnit_5.IN.t12 VGND 0.048675f
C763 distortionUnit_5.IN.n22 VGND 0.084432f
C764 distortionUnit_5.IN.n23 VGND 1.41753f
C765 ui_in[3].t8 VGND 0.01219f
C766 ui_in[3].t18 VGND 0.007184f
C767 ui_in[3].t12 VGND 0.01219f
C768 ui_in[3].t2 VGND 0.007184f
C769 ui_in[3].n0 VGND 0.01758f
C770 ui_in[3].t16 VGND 0.01219f
C771 ui_in[3].t6 VGND 0.007184f
C772 ui_in[3].t15 VGND 0.01219f
C773 ui_in[3].t5 VGND 0.007184f
C774 ui_in[3].n1 VGND 0.01758f
C775 ui_in[3].t17 VGND 0.01219f
C776 ui_in[3].t7 VGND 0.007184f
C777 ui_in[3].n2 VGND 0.016431f
C778 ui_in[3].n3 VGND 0.008046f
C779 ui_in[3].n4 VGND 0.006676f
C780 ui_in[3].n5 VGND 0.008046f
C781 ui_in[3].n6 VGND 0.01758f
C782 ui_in[3].n7 VGND 0.008046f
C783 ui_in[3].n8 VGND 0.006676f
C784 ui_in[3].n9 VGND 0.006676f
C785 ui_in[3].n10 VGND 0.008046f
C786 ui_in[3].n11 VGND 0.01758f
C787 ui_in[3].t9 VGND 0.01219f
C788 ui_in[3].t19 VGND 0.007184f
C789 ui_in[3].t11 VGND 0.01219f
C790 ui_in[3].t1 VGND 0.007184f
C791 ui_in[3].n12 VGND 0.01758f
C792 ui_in[3].t13 VGND 0.01219f
C793 ui_in[3].t3 VGND 0.007184f
C794 ui_in[3].n13 VGND 0.016431f
C795 ui_in[3].n14 VGND 0.008596f
C796 ui_in[3].n15 VGND 0.006676f
C797 ui_in[3].n16 VGND 0.008046f
C798 ui_in[3].n17 VGND 0.01758f
C799 ui_in[3].n18 VGND 0.008046f
C800 ui_in[3].n19 VGND 0.006023f
C801 ui_in[3].n20 VGND 0.409367f
C802 ui_in[3].t14 VGND 0.132645f
C803 ui_in[3].t4 VGND 0.132643f
C804 ui_in[3].n21 VGND 0.767714f
C805 ui_in[3].n22 VGND 0.503797f
C806 ui_in[3].n23 VGND 2.67741f
C807 ui_in[3].t0 VGND 0.136204f
C808 ui_in[3].t10 VGND 0.136202f
C809 ui_in[3].n24 VGND 0.751592f
C810 ui_in[3].n25 VGND 0.509363f
C811 ui_in[3].n26 VGND 1.41582f
C812 ui_in[6].t5 VGND 0.013589f
C813 ui_in[6].t15 VGND 0.008008f
C814 ui_in[6].t7 VGND 0.013589f
C815 ui_in[6].t17 VGND 0.008008f
C816 ui_in[6].n0 VGND 0.019597f
C817 ui_in[6].t6 VGND 0.013589f
C818 ui_in[6].t16 VGND 0.008008f
C819 ui_in[6].t4 VGND 0.013589f
C820 ui_in[6].t14 VGND 0.008008f
C821 ui_in[6].n1 VGND 0.019597f
C822 ui_in[6].t1 VGND 0.013589f
C823 ui_in[6].t12 VGND 0.008008f
C824 ui_in[6].n2 VGND 0.018316f
C825 ui_in[6].n3 VGND 0.008969f
C826 ui_in[6].n4 VGND 0.007442f
C827 ui_in[6].n5 VGND 0.008969f
C828 ui_in[6].n6 VGND 0.019597f
C829 ui_in[6].n7 VGND 0.008969f
C830 ui_in[6].n8 VGND 0.007442f
C831 ui_in[6].n9 VGND 0.007442f
C832 ui_in[6].n10 VGND 0.008969f
C833 ui_in[6].n11 VGND 0.019597f
C834 ui_in[6].t0 VGND 0.013589f
C835 ui_in[6].t11 VGND 0.008008f
C836 ui_in[6].t2 VGND 0.013589f
C837 ui_in[6].t13 VGND 0.008008f
C838 ui_in[6].n12 VGND 0.019597f
C839 ui_in[6].t18 VGND 0.013589f
C840 ui_in[6].t9 VGND 0.008008f
C841 ui_in[6].n13 VGND 0.018316f
C842 ui_in[6].n14 VGND 0.009583f
C843 ui_in[6].n15 VGND 0.007442f
C844 ui_in[6].n16 VGND 0.008969f
C845 ui_in[6].n17 VGND 0.019597f
C846 ui_in[6].n18 VGND 0.008969f
C847 ui_in[6].n19 VGND 0.006714f
C848 ui_in[6].n20 VGND 0.456338f
C849 ui_in[6].t8 VGND 0.147865f
C850 ui_in[6].t10 VGND 0.147863f
C851 ui_in[6].n21 VGND 0.855802f
C852 ui_in[6].n22 VGND 0.561603f
C853 ui_in[6].n23 VGND 2.98462f
C854 ui_in[6].t19 VGND 0.151832f
C855 ui_in[6].t3 VGND 0.15183f
C856 ui_in[6].n24 VGND 0.837831f
C857 ui_in[6].n25 VGND 0.567808f
C858 ui_in[6].n26 VGND 1.57828f
C859 VPWR.n0 VGND 0.624707f
C860 VPWR.n1 VGND 0.67635f
C861 VPWR.n2 VGND 0.110768f
C862 VPWR.n3 VGND 0.110713f
C863 VPWR.n4 VGND 0.221562f
C864 VPWR.n5 VGND 0.221726f
C865 VPWR.n6 VGND 0.673418f
C866 VPWR.n7 VGND 0.110658f
C867 VPWR.n8 VGND 0.111014f
C868 VPWR.n9 VGND 0.661726f
C869 VPWR.n10 VGND 0.110363f
C870 VPWR.n11 VGND 0.110011f
C871 VPWR.n12 VGND 0.220238f
C872 VPWR.n13 VGND 0.660872f
C873 VPWR.n14 VGND 0.675931f
C874 VPWR.n15 VGND 0.66258f
C875 VPWR.n16 VGND 0.220458f
C876 VPWR.n17 VGND 0.110201f
C877 VPWR.n18 VGND 0.110255f
C878 VPWR.n19 VGND 0.379109f
C879 VPWR.n20 VGND 0.707327f
C880 VPWR.t265 VGND 0.038813f
C881 VPWR.t267 VGND 0.00879f
C882 VPWR.n21 VGND 0.05086f
C883 VPWR.t74 VGND 0.002392f
C884 VPWR.t58 VGND 0.002392f
C885 VPWR.n22 VGND 0.004947f
C886 VPWR.n23 VGND 0.098234f
C887 VPWR.t62 VGND 0.002392f
C888 VPWR.t66 VGND 0.002392f
C889 VPWR.n24 VGND 0.004947f
C890 VPWR.n25 VGND 0.082582f
C891 VPWR.t259 VGND 0.038787f
C892 VPWR.t261 VGND 0.00879f
C893 VPWR.n26 VGND 0.090806f
C894 VPWR.t64 VGND 0.002392f
C895 VPWR.t68 VGND 0.002392f
C896 VPWR.n27 VGND 0.004947f
C897 VPWR.n28 VGND 0.119761f
C898 VPWR.t76 VGND 0.002392f
C899 VPWR.t60 VGND 0.002392f
C900 VPWR.n29 VGND 0.004947f
C901 VPWR.n30 VGND 0.072188f
C902 VPWR.t266 VGND 0.136425f
C903 VPWR.t73 VGND 0.108971f
C904 VPWR.t57 VGND 0.108971f
C905 VPWR.t61 VGND 0.108971f
C906 VPWR.t65 VGND 0.108971f
C907 VPWR.t69 VGND 0.078349f
C908 VPWR.t260 VGND 0.136425f
C909 VPWR.t67 VGND 0.108971f
C910 VPWR.t63 VGND 0.108971f
C911 VPWR.t59 VGND 0.108971f
C912 VPWR.t75 VGND 0.108971f
C913 VPWR.t71 VGND 0.085107f
C914 VPWR.n31 VGND -0.063904f
C915 VPWR.t107 VGND 0.091784f
C916 VPWR.n32 VGND 0.140992f
C917 VPWR.n33 VGND 0.018809f
C918 VPWR.t70 VGND 0.002392f
C919 VPWR.t72 VGND 0.002392f
C920 VPWR.n34 VGND 0.004947f
C921 VPWR.n35 VGND 0.081171f
C922 VPWR.n36 VGND 2.89145f
C923 VPWR.n37 VGND 1.42069f
C924 VPWR.n38 VGND 0.003801f
C925 VPWR.n39 VGND 0.007286f
C926 VPWR.t47 VGND 0.002227f
C927 VPWR.t11 VGND 0.002227f
C928 VPWR.n40 VGND 0.004781f
C929 VPWR.t12 VGND 0.002227f
C930 VPWR.t110 VGND 0.002227f
C931 VPWR.n41 VGND 0.004781f
C932 VPWR.n42 VGND 0.001991f
C933 VPWR.t111 VGND 0.00848f
C934 VPWR.n43 VGND 0.012082f
C935 VPWR.n44 VGND 0.005464f
C936 VPWR.n45 VGND 0.007286f
C937 VPWR.n46 VGND 0.007286f
C938 VPWR.n47 VGND 0.001416f
C939 VPWR.n48 VGND 0.005451f
C940 VPWR.n49 VGND 0.002356f
C941 VPWR.n50 VGND 0.005451f
C942 VPWR.t109 VGND 0.002227f
C943 VPWR.t10 VGND 0.002227f
C944 VPWR.n51 VGND 0.004781f
C945 VPWR.n52 VGND 0.001795f
C946 VPWR.t48 VGND 0.008481f
C947 VPWR.n53 VGND 0.009967f
C948 VPWR.n54 VGND 0.004545f
C949 VPWR.n55 VGND 0.007286f
C950 VPWR.n56 VGND 0.007286f
C951 VPWR.n57 VGND 0.001613f
C952 VPWR.n58 VGND 0.005451f
C953 VPWR.n59 VGND 0.002258f
C954 VPWR.n60 VGND 0.001388f
C955 VPWR.n61 VGND 0.007127f
C956 VPWR.n62 VGND 0.292827f
C957 VPWR.n63 VGND 0.029122f
C958 VPWR.n64 VGND 0.016784f
C959 VPWR.n65 VGND 0.119794f
C960 VPWR.t46 VGND 0.095507f
C961 VPWR.n66 VGND 0.060445f
C962 VPWR.t287 VGND 0.095507f
C963 VPWR.n67 VGND 0.098959f
C964 VPWR.n68 VGND 0.05179f
C965 VPWR.n69 VGND 0.228182f
C966 VPWR.n70 VGND 0.029122f
C967 VPWR.n71 VGND 0.016784f
C968 VPWR.n72 VGND 0.119794f
C969 VPWR.t97 VGND 0.095507f
C970 VPWR.n73 VGND 0.060445f
C971 VPWR.t98 VGND 0.095507f
C972 VPWR.n74 VGND 0.098959f
C973 VPWR.n75 VGND 0.05179f
C974 VPWR.n76 VGND 0.23101f
C975 VPWR.n77 VGND 0.212637f
C976 VPWR.n78 VGND 29.132902f
C977 VPWR.n79 VGND 0.624707f
C978 VPWR.n80 VGND 0.67635f
C979 VPWR.n81 VGND 0.110768f
C980 VPWR.n82 VGND 0.110713f
C981 VPWR.n83 VGND 0.221562f
C982 VPWR.n84 VGND 0.221726f
C983 VPWR.n85 VGND 0.673418f
C984 VPWR.n86 VGND 0.110658f
C985 VPWR.n87 VGND 0.111014f
C986 VPWR.n88 VGND 0.661726f
C987 VPWR.n89 VGND 0.110363f
C988 VPWR.n90 VGND 0.110011f
C989 VPWR.n91 VGND 0.220238f
C990 VPWR.n92 VGND 0.660872f
C991 VPWR.n93 VGND 0.675931f
C992 VPWR.n94 VGND 0.66258f
C993 VPWR.n95 VGND 0.220458f
C994 VPWR.n96 VGND 0.110201f
C995 VPWR.n97 VGND 0.110255f
C996 VPWR.n98 VGND 0.379109f
C997 VPWR.n99 VGND 0.707327f
C998 VPWR.t250 VGND 0.038813f
C999 VPWR.t252 VGND 0.00879f
C1000 VPWR.n100 VGND 0.05086f
C1001 VPWR.t213 VGND 0.002392f
C1002 VPWR.t223 VGND 0.002392f
C1003 VPWR.n101 VGND 0.004947f
C1004 VPWR.n102 VGND 0.098234f
C1005 VPWR.t227 VGND 0.002392f
C1006 VPWR.t211 VGND 0.002392f
C1007 VPWR.n103 VGND 0.004947f
C1008 VPWR.n104 VGND 0.082582f
C1009 VPWR.t244 VGND 0.038787f
C1010 VPWR.t246 VGND 0.00879f
C1011 VPWR.n105 VGND 0.090806f
C1012 VPWR.t209 VGND 0.002392f
C1013 VPWR.t215 VGND 0.002392f
C1014 VPWR.n106 VGND 0.004947f
C1015 VPWR.n107 VGND 0.119761f
C1016 VPWR.t221 VGND 0.002392f
C1017 VPWR.t225 VGND 0.002392f
C1018 VPWR.n108 VGND 0.004947f
C1019 VPWR.n109 VGND 0.072188f
C1020 VPWR.t251 VGND 0.136425f
C1021 VPWR.t212 VGND 0.108971f
C1022 VPWR.t222 VGND 0.108971f
C1023 VPWR.t226 VGND 0.108971f
C1024 VPWR.t210 VGND 0.108971f
C1025 VPWR.t218 VGND 0.078349f
C1026 VPWR.t245 VGND 0.136425f
C1027 VPWR.t214 VGND 0.108971f
C1028 VPWR.t208 VGND 0.108971f
C1029 VPWR.t224 VGND 0.108971f
C1030 VPWR.t220 VGND 0.108971f
C1031 VPWR.t216 VGND 0.085107f
C1032 VPWR.n110 VGND -0.063904f
C1033 VPWR.t106 VGND 0.091784f
C1034 VPWR.n111 VGND 0.140992f
C1035 VPWR.n112 VGND 0.018809f
C1036 VPWR.t219 VGND 0.002392f
C1037 VPWR.t217 VGND 0.002392f
C1038 VPWR.n113 VGND 0.004947f
C1039 VPWR.n114 VGND 0.081171f
C1040 VPWR.n115 VGND 2.89145f
C1041 VPWR.n116 VGND 1.42069f
C1042 VPWR.n117 VGND 0.003801f
C1043 VPWR.n118 VGND 0.007286f
C1044 VPWR.t103 VGND 0.002227f
C1045 VPWR.t228 VGND 0.002227f
C1046 VPWR.n119 VGND 0.004781f
C1047 VPWR.t50 VGND 0.002227f
C1048 VPWR.t87 VGND 0.002227f
C1049 VPWR.n120 VGND 0.004781f
C1050 VPWR.n121 VGND 0.001991f
C1051 VPWR.t104 VGND 0.00848f
C1052 VPWR.n122 VGND 0.012082f
C1053 VPWR.n123 VGND 0.005464f
C1054 VPWR.n124 VGND 0.007286f
C1055 VPWR.n125 VGND 0.007286f
C1056 VPWR.n126 VGND 0.001416f
C1057 VPWR.n127 VGND 0.005451f
C1058 VPWR.n128 VGND 0.002356f
C1059 VPWR.n129 VGND 0.005451f
C1060 VPWR.t89 VGND 0.002227f
C1061 VPWR.t49 VGND 0.002227f
C1062 VPWR.n130 VGND 0.004781f
C1063 VPWR.n131 VGND 0.001795f
C1064 VPWR.t86 VGND 0.008481f
C1065 VPWR.n132 VGND 0.009967f
C1066 VPWR.n133 VGND 0.004545f
C1067 VPWR.n134 VGND 0.007286f
C1068 VPWR.n135 VGND 0.007286f
C1069 VPWR.n136 VGND 0.001613f
C1070 VPWR.n137 VGND 0.005451f
C1071 VPWR.n138 VGND 0.002258f
C1072 VPWR.n139 VGND 0.001388f
C1073 VPWR.n140 VGND 0.007127f
C1074 VPWR.n141 VGND 0.292827f
C1075 VPWR.n142 VGND 0.029122f
C1076 VPWR.n143 VGND 0.016784f
C1077 VPWR.n144 VGND 0.119794f
C1078 VPWR.t105 VGND 0.095507f
C1079 VPWR.n145 VGND 0.060445f
C1080 VPWR.t88 VGND 0.095507f
C1081 VPWR.n146 VGND 0.098959f
C1082 VPWR.n147 VGND 0.05179f
C1083 VPWR.n148 VGND 0.228182f
C1084 VPWR.n149 VGND 0.029122f
C1085 VPWR.n150 VGND 0.016784f
C1086 VPWR.n151 VGND 0.119794f
C1087 VPWR.t78 VGND 0.095507f
C1088 VPWR.n152 VGND 0.060445f
C1089 VPWR.t79 VGND 0.095507f
C1090 VPWR.n153 VGND 0.098959f
C1091 VPWR.n154 VGND 0.05179f
C1092 VPWR.n155 VGND 0.23101f
C1093 VPWR.n156 VGND 0.212637f
C1094 VPWR.n157 VGND 5.0391f
C1095 VPWR.n158 VGND 0.415614p
C1096 VPWR.n159 VGND 15.439699f
C1097 VPWR.n160 VGND 0.624707f
C1098 VPWR.n161 VGND 0.67635f
C1099 VPWR.n162 VGND 0.110768f
C1100 VPWR.n163 VGND 0.110713f
C1101 VPWR.n164 VGND 0.221562f
C1102 VPWR.n165 VGND 0.221726f
C1103 VPWR.n166 VGND 0.673418f
C1104 VPWR.n167 VGND 0.110658f
C1105 VPWR.n168 VGND 0.111014f
C1106 VPWR.n169 VGND 0.661726f
C1107 VPWR.n170 VGND 0.110363f
C1108 VPWR.n171 VGND 0.110011f
C1109 VPWR.n172 VGND 0.220238f
C1110 VPWR.n173 VGND 0.660872f
C1111 VPWR.n174 VGND 0.675931f
C1112 VPWR.n175 VGND 0.66258f
C1113 VPWR.n176 VGND 0.220458f
C1114 VPWR.n177 VGND 0.110201f
C1115 VPWR.n178 VGND 0.110255f
C1116 VPWR.n179 VGND 0.379109f
C1117 VPWR.n180 VGND 0.707327f
C1118 VPWR.t253 VGND 0.038813f
C1119 VPWR.t255 VGND 0.00879f
C1120 VPWR.n181 VGND 0.05086f
C1121 VPWR.t299 VGND 0.002392f
C1122 VPWR.t305 VGND 0.002392f
C1123 VPWR.n182 VGND 0.004947f
C1124 VPWR.n183 VGND 0.098234f
C1125 VPWR.t309 VGND 0.002392f
C1126 VPWR.t297 VGND 0.002392f
C1127 VPWR.n184 VGND 0.004947f
C1128 VPWR.n185 VGND 0.082582f
C1129 VPWR.t247 VGND 0.038787f
C1130 VPWR.t249 VGND 0.00879f
C1131 VPWR.n186 VGND 0.090806f
C1132 VPWR.t293 VGND 0.002392f
C1133 VPWR.t311 VGND 0.002392f
C1134 VPWR.n187 VGND 0.004947f
C1135 VPWR.n188 VGND 0.119761f
C1136 VPWR.t303 VGND 0.002392f
C1137 VPWR.t307 VGND 0.002392f
C1138 VPWR.n189 VGND 0.004947f
C1139 VPWR.n190 VGND 0.072188f
C1140 VPWR.t254 VGND 0.136425f
C1141 VPWR.t298 VGND 0.108971f
C1142 VPWR.t304 VGND 0.108971f
C1143 VPWR.t308 VGND 0.108971f
C1144 VPWR.t296 VGND 0.108971f
C1145 VPWR.t294 VGND 0.078349f
C1146 VPWR.t248 VGND 0.136425f
C1147 VPWR.t310 VGND 0.108971f
C1148 VPWR.t292 VGND 0.108971f
C1149 VPWR.t306 VGND 0.108971f
C1150 VPWR.t302 VGND 0.108971f
C1151 VPWR.t300 VGND 0.085107f
C1152 VPWR.n191 VGND -0.063904f
C1153 VPWR.t95 VGND 0.091784f
C1154 VPWR.n192 VGND 0.140992f
C1155 VPWR.n193 VGND 0.018809f
C1156 VPWR.t295 VGND 0.002392f
C1157 VPWR.t301 VGND 0.002392f
C1158 VPWR.n194 VGND 0.004947f
C1159 VPWR.n195 VGND 0.081171f
C1160 VPWR.n196 VGND 2.89145f
C1161 VPWR.n197 VGND 1.42069f
C1162 VPWR.n198 VGND 0.003801f
C1163 VPWR.n199 VGND 0.007286f
C1164 VPWR.t80 VGND 0.002227f
C1165 VPWR.t33 VGND 0.002227f
C1166 VPWR.n200 VGND 0.004781f
C1167 VPWR.t100 VGND 0.002227f
C1168 VPWR.t34 VGND 0.002227f
C1169 VPWR.n201 VGND 0.004781f
C1170 VPWR.n202 VGND 0.001991f
C1171 VPWR.t81 VGND 0.00848f
C1172 VPWR.n203 VGND 0.012082f
C1173 VPWR.n204 VGND 0.005464f
C1174 VPWR.n205 VGND 0.007286f
C1175 VPWR.n206 VGND 0.007286f
C1176 VPWR.n207 VGND 0.001416f
C1177 VPWR.n208 VGND 0.005451f
C1178 VPWR.n209 VGND 0.002356f
C1179 VPWR.n210 VGND 0.005451f
C1180 VPWR.t102 VGND 0.002227f
C1181 VPWR.t99 VGND 0.002227f
C1182 VPWR.n211 VGND 0.004781f
C1183 VPWR.n212 VGND 0.001795f
C1184 VPWR.t101 VGND 0.008481f
C1185 VPWR.n213 VGND 0.009967f
C1186 VPWR.n214 VGND 0.004545f
C1187 VPWR.n215 VGND 0.007286f
C1188 VPWR.n216 VGND 0.007286f
C1189 VPWR.n217 VGND 0.001613f
C1190 VPWR.n218 VGND 0.005451f
C1191 VPWR.n219 VGND 0.002258f
C1192 VPWR.n220 VGND 0.001388f
C1193 VPWR.n221 VGND 0.007127f
C1194 VPWR.n222 VGND 0.292827f
C1195 VPWR.n223 VGND 0.029122f
C1196 VPWR.n224 VGND 0.016784f
C1197 VPWR.n225 VGND 0.119794f
C1198 VPWR.t35 VGND 0.095507f
C1199 VPWR.n226 VGND 0.060445f
C1200 VPWR.t54 VGND 0.095507f
C1201 VPWR.n227 VGND 0.098959f
C1202 VPWR.n228 VGND 0.05179f
C1203 VPWR.n229 VGND 0.228182f
C1204 VPWR.n230 VGND 0.029122f
C1205 VPWR.n231 VGND 0.016784f
C1206 VPWR.n232 VGND 0.119794f
C1207 VPWR.t279 VGND 0.095507f
C1208 VPWR.n233 VGND 0.060445f
C1209 VPWR.t280 VGND 0.095507f
C1210 VPWR.n234 VGND 0.098959f
C1211 VPWR.n235 VGND 0.05179f
C1212 VPWR.n236 VGND 0.23101f
C1213 VPWR.n237 VGND 0.212637f
C1214 VPWR.n238 VGND 12.653f
C1215 VPWR.n239 VGND 0.624707f
C1216 VPWR.n240 VGND 0.67635f
C1217 VPWR.n241 VGND 0.110768f
C1218 VPWR.n242 VGND 0.110713f
C1219 VPWR.n243 VGND 0.221562f
C1220 VPWR.n244 VGND 0.221726f
C1221 VPWR.n245 VGND 0.673418f
C1222 VPWR.n246 VGND 0.110658f
C1223 VPWR.n247 VGND 0.111014f
C1224 VPWR.n248 VGND 0.661726f
C1225 VPWR.n249 VGND 0.110363f
C1226 VPWR.n250 VGND 0.110011f
C1227 VPWR.n251 VGND 0.220238f
C1228 VPWR.n252 VGND 0.660872f
C1229 VPWR.n253 VGND 0.675931f
C1230 VPWR.n254 VGND 0.66258f
C1231 VPWR.n255 VGND 0.220458f
C1232 VPWR.n256 VGND 0.110201f
C1233 VPWR.n257 VGND 0.110255f
C1234 VPWR.n258 VGND 0.379109f
C1235 VPWR.n259 VGND 0.707327f
C1236 VPWR.t235 VGND 0.038813f
C1237 VPWR.t237 VGND 0.00879f
C1238 VPWR.n260 VGND 0.05086f
C1239 VPWR.t142 VGND 0.002392f
C1240 VPWR.t146 VGND 0.002392f
C1241 VPWR.n261 VGND 0.004947f
C1242 VPWR.n262 VGND 0.098234f
C1243 VPWR.t152 VGND 0.002392f
C1244 VPWR.t138 VGND 0.002392f
C1245 VPWR.n263 VGND 0.004947f
C1246 VPWR.n264 VGND 0.082582f
C1247 VPWR.t241 VGND 0.038787f
C1248 VPWR.t243 VGND 0.00879f
C1249 VPWR.n265 VGND 0.090806f
C1250 VPWR.t148 VGND 0.002392f
C1251 VPWR.t154 VGND 0.002392f
C1252 VPWR.n266 VGND 0.004947f
C1253 VPWR.n267 VGND 0.119761f
C1254 VPWR.t144 VGND 0.002392f
C1255 VPWR.t150 VGND 0.002392f
C1256 VPWR.n268 VGND 0.004947f
C1257 VPWR.n269 VGND 0.072188f
C1258 VPWR.t236 VGND 0.136425f
C1259 VPWR.t141 VGND 0.108971f
C1260 VPWR.t145 VGND 0.108971f
C1261 VPWR.t151 VGND 0.108971f
C1262 VPWR.t137 VGND 0.108971f
C1263 VPWR.t155 VGND 0.078349f
C1264 VPWR.t242 VGND 0.136425f
C1265 VPWR.t153 VGND 0.108971f
C1266 VPWR.t147 VGND 0.108971f
C1267 VPWR.t149 VGND 0.108971f
C1268 VPWR.t143 VGND 0.108971f
C1269 VPWR.t139 VGND 0.085107f
C1270 VPWR.n270 VGND -0.063904f
C1271 VPWR.t108 VGND 0.091784f
C1272 VPWR.n271 VGND 0.140992f
C1273 VPWR.n272 VGND 0.018809f
C1274 VPWR.t156 VGND 0.002392f
C1275 VPWR.t140 VGND 0.002392f
C1276 VPWR.n273 VGND 0.004947f
C1277 VPWR.n274 VGND 0.081171f
C1278 VPWR.n275 VGND 2.89145f
C1279 VPWR.n276 VGND 1.42069f
C1280 VPWR.n277 VGND 0.003801f
C1281 VPWR.n278 VGND 0.007286f
C1282 VPWR.t160 VGND 0.002227f
C1283 VPWR.t96 VGND 0.002227f
C1284 VPWR.n279 VGND 0.004781f
C1285 VPWR.t36 VGND 0.002227f
C1286 VPWR.t37 VGND 0.002227f
C1287 VPWR.n280 VGND 0.004781f
C1288 VPWR.n281 VGND 0.001991f
C1289 VPWR.t38 VGND 0.00848f
C1290 VPWR.n282 VGND 0.012082f
C1291 VPWR.n283 VGND 0.005464f
C1292 VPWR.n284 VGND 0.007286f
C1293 VPWR.n285 VGND 0.007286f
C1294 VPWR.n286 VGND 0.001416f
C1295 VPWR.n287 VGND 0.005451f
C1296 VPWR.n288 VGND 0.002356f
C1297 VPWR.n289 VGND 0.005451f
C1298 VPWR.t157 VGND 0.002227f
C1299 VPWR.t159 VGND 0.002227f
C1300 VPWR.n290 VGND 0.004781f
C1301 VPWR.n291 VGND 0.001795f
C1302 VPWR.t161 VGND 0.008481f
C1303 VPWR.n292 VGND 0.009967f
C1304 VPWR.n293 VGND 0.004545f
C1305 VPWR.n294 VGND 0.007286f
C1306 VPWR.n295 VGND 0.007286f
C1307 VPWR.n296 VGND 0.001613f
C1308 VPWR.n297 VGND 0.005451f
C1309 VPWR.n298 VGND 0.002258f
C1310 VPWR.n299 VGND 0.001388f
C1311 VPWR.n300 VGND 0.007127f
C1312 VPWR.n301 VGND 0.292827f
C1313 VPWR.n302 VGND 0.029122f
C1314 VPWR.n303 VGND 0.016784f
C1315 VPWR.n304 VGND 0.119794f
C1316 VPWR.t158 VGND 0.095507f
C1317 VPWR.n305 VGND 0.060445f
C1318 VPWR.t278 VGND 0.095507f
C1319 VPWR.n306 VGND 0.098959f
C1320 VPWR.n307 VGND 0.05179f
C1321 VPWR.n308 VGND 0.228182f
C1322 VPWR.n309 VGND 0.029122f
C1323 VPWR.n310 VGND 0.016784f
C1324 VPWR.n311 VGND 0.119794f
C1325 VPWR.t206 VGND 0.095507f
C1326 VPWR.n312 VGND 0.060445f
C1327 VPWR.t207 VGND 0.095507f
C1328 VPWR.n313 VGND 0.098959f
C1329 VPWR.n314 VGND 0.05179f
C1330 VPWR.n315 VGND 0.23101f
C1331 VPWR.n316 VGND 0.212637f
C1332 VPWR.n317 VGND 5.0391f
C1333 VPWR.n318 VGND 0.346915p
C1334 VPWR.n319 VGND 0.029122f
C1335 VPWR.n320 VGND 0.016784f
C1336 VPWR.n321 VGND 0.119794f
C1337 VPWR.t289 VGND 0.095507f
C1338 VPWR.n322 VGND 0.060445f
C1339 VPWR.t134 VGND 0.095507f
C1340 VPWR.n323 VGND 0.098959f
C1341 VPWR.n324 VGND 0.05179f
C1342 VPWR.n325 VGND 0.228182f
C1343 VPWR.n326 VGND 0.029122f
C1344 VPWR.n327 VGND 0.016784f
C1345 VPWR.n328 VGND 0.119794f
C1346 VPWR.t55 VGND 0.095507f
C1347 VPWR.n329 VGND 0.060445f
C1348 VPWR.t56 VGND 0.095507f
C1349 VPWR.n330 VGND 0.098959f
C1350 VPWR.n331 VGND 0.05179f
C1351 VPWR.n332 VGND 0.23101f
C1352 VPWR.n333 VGND 0.512436f
C1353 VPWR.n334 VGND 0.003801f
C1354 VPWR.n335 VGND 0.007286f
C1355 VPWR.t290 VGND 0.002227f
C1356 VPWR.t133 VGND 0.002227f
C1357 VPWR.n336 VGND 0.004781f
C1358 VPWR.t112 VGND 0.002227f
C1359 VPWR.t135 VGND 0.002227f
C1360 VPWR.n337 VGND 0.004781f
C1361 VPWR.n338 VGND 0.001991f
C1362 VPWR.t136 VGND 0.00848f
C1363 VPWR.n339 VGND 0.012082f
C1364 VPWR.n340 VGND 0.005464f
C1365 VPWR.n341 VGND 0.007286f
C1366 VPWR.n342 VGND 0.007286f
C1367 VPWR.n343 VGND 0.001416f
C1368 VPWR.n344 VGND 0.005451f
C1369 VPWR.n345 VGND 0.002356f
C1370 VPWR.n346 VGND 0.005451f
C1371 VPWR.t185 VGND 0.002227f
C1372 VPWR.t288 VGND 0.002227f
C1373 VPWR.n347 VGND 0.004781f
C1374 VPWR.n348 VGND 0.001795f
C1375 VPWR.t291 VGND 0.008481f
C1376 VPWR.n349 VGND 0.009967f
C1377 VPWR.n350 VGND 0.004545f
C1378 VPWR.n351 VGND 0.007286f
C1379 VPWR.n352 VGND 0.007286f
C1380 VPWR.n353 VGND 0.001613f
C1381 VPWR.n354 VGND 0.005451f
C1382 VPWR.n355 VGND 0.002258f
C1383 VPWR.n356 VGND 0.001388f
C1384 VPWR.n357 VGND 0.007127f
C1385 VPWR.n358 VGND 0.292827f
C1386 VPWR.n359 VGND 7.28225f
C1387 VPWR.n360 VGND 0.624707f
C1388 VPWR.n361 VGND 0.67635f
C1389 VPWR.n362 VGND 0.110768f
C1390 VPWR.n363 VGND 0.110713f
C1391 VPWR.n364 VGND 0.221562f
C1392 VPWR.n365 VGND 0.221726f
C1393 VPWR.n366 VGND 0.673418f
C1394 VPWR.n367 VGND 0.110658f
C1395 VPWR.n368 VGND 0.111014f
C1396 VPWR.n369 VGND 0.661726f
C1397 VPWR.n370 VGND 0.110363f
C1398 VPWR.n371 VGND 0.110011f
C1399 VPWR.n372 VGND 0.220238f
C1400 VPWR.n373 VGND 0.660872f
C1401 VPWR.n374 VGND 0.675931f
C1402 VPWR.n375 VGND 0.66258f
C1403 VPWR.n376 VGND 0.220458f
C1404 VPWR.n377 VGND 0.110201f
C1405 VPWR.n378 VGND 0.110255f
C1406 VPWR.n379 VGND 0.379109f
C1407 VPWR.n380 VGND 0.707327f
C1408 VPWR.t232 VGND 0.038813f
C1409 VPWR.t234 VGND 0.00879f
C1410 VPWR.n381 VGND 0.05086f
C1411 VPWR.t195 VGND 0.002392f
C1412 VPWR.t193 VGND 0.002392f
C1413 VPWR.n382 VGND 0.004947f
C1414 VPWR.n383 VGND 0.098234f
C1415 VPWR.t199 VGND 0.002392f
C1416 VPWR.t187 VGND 0.002392f
C1417 VPWR.n384 VGND 0.004947f
C1418 VPWR.n385 VGND 0.082582f
C1419 VPWR.t238 VGND 0.038787f
C1420 VPWR.t240 VGND 0.00879f
C1421 VPWR.n386 VGND 0.090806f
C1422 VPWR.t201 VGND 0.002392f
C1423 VPWR.t203 VGND 0.002392f
C1424 VPWR.n387 VGND 0.004947f
C1425 VPWR.n388 VGND 0.119761f
C1426 VPWR.t189 VGND 0.002392f
C1427 VPWR.t197 VGND 0.002392f
C1428 VPWR.n389 VGND 0.004947f
C1429 VPWR.n390 VGND 0.072188f
C1430 VPWR.t233 VGND 0.136425f
C1431 VPWR.t194 VGND 0.108971f
C1432 VPWR.t192 VGND 0.108971f
C1433 VPWR.t198 VGND 0.108971f
C1434 VPWR.t186 VGND 0.108971f
C1435 VPWR.t204 VGND 0.078349f
C1436 VPWR.t239 VGND 0.136425f
C1437 VPWR.t202 VGND 0.108971f
C1438 VPWR.t200 VGND 0.108971f
C1439 VPWR.t196 VGND 0.108971f
C1440 VPWR.t188 VGND 0.108971f
C1441 VPWR.t190 VGND 0.085107f
C1442 VPWR.n391 VGND -0.063904f
C1443 VPWR.t277 VGND 0.091784f
C1444 VPWR.n392 VGND 0.140992f
C1445 VPWR.n393 VGND 0.018809f
C1446 VPWR.t205 VGND 0.002392f
C1447 VPWR.t191 VGND 0.002392f
C1448 VPWR.n394 VGND 0.004947f
C1449 VPWR.n395 VGND 0.081171f
C1450 VPWR.n396 VGND 2.89145f
C1451 VPWR.n397 VGND 1.42069f
C1452 VPWR.n398 VGND 4.94303f
C1453 VPWR.n399 VGND 0.029122f
C1454 VPWR.n400 VGND 0.016784f
C1455 VPWR.n401 VGND 0.119794f
C1456 VPWR.t8 VGND 0.095507f
C1457 VPWR.n402 VGND 0.060445f
C1458 VPWR.t0 VGND 0.095507f
C1459 VPWR.n403 VGND 0.098959f
C1460 VPWR.n404 VGND 0.05179f
C1461 VPWR.n405 VGND 0.228182f
C1462 VPWR.n406 VGND 0.029122f
C1463 VPWR.n407 VGND 0.016784f
C1464 VPWR.n408 VGND 0.119794f
C1465 VPWR.t53 VGND 0.095507f
C1466 VPWR.n409 VGND 0.060445f
C1467 VPWR.t52 VGND 0.095507f
C1468 VPWR.n410 VGND 0.098959f
C1469 VPWR.n411 VGND 0.05179f
C1470 VPWR.n412 VGND 0.23101f
C1471 VPWR.n413 VGND 0.212637f
C1472 VPWR.n414 VGND 3.44362f
C1473 VPWR.n415 VGND 0.003801f
C1474 VPWR.n416 VGND 0.007286f
C1475 VPWR.t6 VGND 0.002227f
C1476 VPWR.t4 VGND 0.002227f
C1477 VPWR.n417 VGND 0.004781f
C1478 VPWR.t3 VGND 0.002227f
C1479 VPWR.t1 VGND 0.002227f
C1480 VPWR.n418 VGND 0.004781f
C1481 VPWR.n419 VGND 0.001991f
C1482 VPWR.t5 VGND 0.00848f
C1483 VPWR.n420 VGND 0.012082f
C1484 VPWR.n421 VGND 0.005464f
C1485 VPWR.n422 VGND 0.007286f
C1486 VPWR.n423 VGND 0.007286f
C1487 VPWR.n424 VGND 0.001416f
C1488 VPWR.n425 VGND 0.005451f
C1489 VPWR.n426 VGND 0.002356f
C1490 VPWR.n427 VGND 0.005451f
C1491 VPWR.t7 VGND 0.002227f
C1492 VPWR.t9 VGND 0.002227f
C1493 VPWR.n428 VGND 0.004781f
C1494 VPWR.n429 VGND 0.001795f
C1495 VPWR.t2 VGND 0.008481f
C1496 VPWR.n430 VGND 0.009967f
C1497 VPWR.n431 VGND 0.004545f
C1498 VPWR.n432 VGND 0.007286f
C1499 VPWR.n433 VGND 0.007286f
C1500 VPWR.n434 VGND 0.001613f
C1501 VPWR.n435 VGND 0.005451f
C1502 VPWR.n436 VGND 0.002258f
C1503 VPWR.n437 VGND 0.001388f
C1504 VPWR.n438 VGND 0.007127f
C1505 VPWR.n439 VGND 0.292827f
C1506 VPWR.n440 VGND 4.84854f
C1507 VPWR.n441 VGND 0.624707f
C1508 VPWR.n442 VGND 0.67635f
C1509 VPWR.n443 VGND 0.110768f
C1510 VPWR.n444 VGND 0.110713f
C1511 VPWR.n445 VGND 0.221562f
C1512 VPWR.n446 VGND 0.221726f
C1513 VPWR.n447 VGND 0.673418f
C1514 VPWR.n448 VGND 0.110658f
C1515 VPWR.n449 VGND 0.111014f
C1516 VPWR.n450 VGND 0.661726f
C1517 VPWR.n451 VGND 0.110363f
C1518 VPWR.n452 VGND 0.110011f
C1519 VPWR.n453 VGND 0.220238f
C1520 VPWR.n454 VGND 0.660872f
C1521 VPWR.n455 VGND 0.675931f
C1522 VPWR.n456 VGND 0.66258f
C1523 VPWR.n457 VGND 0.220458f
C1524 VPWR.n458 VGND 0.110201f
C1525 VPWR.n459 VGND 0.110255f
C1526 VPWR.n460 VGND 0.379109f
C1527 VPWR.n461 VGND 0.707327f
C1528 VPWR.t229 VGND 0.038813f
C1529 VPWR.t231 VGND 0.00879f
C1530 VPWR.n462 VGND 0.05086f
C1531 VPWR.t24 VGND 0.002392f
C1532 VPWR.t28 VGND 0.002392f
C1533 VPWR.n463 VGND 0.004947f
C1534 VPWR.n464 VGND 0.098234f
C1535 VPWR.t32 VGND 0.002392f
C1536 VPWR.t20 VGND 0.002392f
C1537 VPWR.n465 VGND 0.004947f
C1538 VPWR.n466 VGND 0.082582f
C1539 VPWR.t256 VGND 0.038787f
C1540 VPWR.t258 VGND 0.00879f
C1541 VPWR.n467 VGND 0.090806f
C1542 VPWR.t16 VGND 0.002392f
C1543 VPWR.t14 VGND 0.002392f
C1544 VPWR.n468 VGND 0.004947f
C1545 VPWR.n469 VGND 0.119761f
C1546 VPWR.t22 VGND 0.002392f
C1547 VPWR.t30 VGND 0.002392f
C1548 VPWR.n470 VGND 0.004947f
C1549 VPWR.n471 VGND 0.072188f
C1550 VPWR.t230 VGND 0.136425f
C1551 VPWR.t23 VGND 0.108971f
C1552 VPWR.t27 VGND 0.108971f
C1553 VPWR.t31 VGND 0.108971f
C1554 VPWR.t19 VGND 0.108971f
C1555 VPWR.t17 VGND 0.078349f
C1556 VPWR.t257 VGND 0.136425f
C1557 VPWR.t13 VGND 0.108971f
C1558 VPWR.t15 VGND 0.108971f
C1559 VPWR.t29 VGND 0.108971f
C1560 VPWR.t21 VGND 0.108971f
C1561 VPWR.t25 VGND 0.085107f
C1562 VPWR.n472 VGND -0.063904f
C1563 VPWR.t51 VGND 0.091784f
C1564 VPWR.n473 VGND 0.140992f
C1565 VPWR.n474 VGND 0.018809f
C1566 VPWR.t18 VGND 0.002392f
C1567 VPWR.t26 VGND 0.002392f
C1568 VPWR.n475 VGND 0.004947f
C1569 VPWR.n476 VGND 0.081171f
C1570 VPWR.n477 VGND 2.89145f
C1571 VPWR.n478 VGND 1.42069f
C1572 VPWR.n479 VGND 4.94303f
C1573 VPWR.n480 VGND 7.5835f
C1574 VPWR.n481 VGND 0.029122f
C1575 VPWR.n482 VGND 0.016784f
C1576 VPWR.n483 VGND 0.119794f
C1577 VPWR.t90 VGND 0.095507f
C1578 VPWR.n484 VGND 0.060445f
C1579 VPWR.t77 VGND 0.095507f
C1580 VPWR.n485 VGND 0.098959f
C1581 VPWR.n486 VGND 0.05179f
C1582 VPWR.n487 VGND 0.228182f
C1583 VPWR.n488 VGND 0.029122f
C1584 VPWR.n489 VGND 0.016784f
C1585 VPWR.n490 VGND 0.119794f
C1586 VPWR.t285 VGND 0.095507f
C1587 VPWR.n491 VGND 0.060445f
C1588 VPWR.t286 VGND 0.095507f
C1589 VPWR.n492 VGND 0.098959f
C1590 VPWR.n493 VGND 0.05179f
C1591 VPWR.n494 VGND 0.23101f
C1592 VPWR.n495 VGND 0.452983f
C1593 VPWR.n496 VGND 0.003801f
C1594 VPWR.n497 VGND 0.007286f
C1595 VPWR.t94 VGND 0.002227f
C1596 VPWR.t84 VGND 0.002227f
C1597 VPWR.n498 VGND 0.004781f
C1598 VPWR.t85 VGND 0.002227f
C1599 VPWR.t93 VGND 0.002227f
C1600 VPWR.n499 VGND 0.004781f
C1601 VPWR.n500 VGND 0.001991f
C1602 VPWR.t82 VGND 0.00848f
C1603 VPWR.n501 VGND 0.012082f
C1604 VPWR.n502 VGND 0.005464f
C1605 VPWR.n503 VGND 0.007286f
C1606 VPWR.n504 VGND 0.007286f
C1607 VPWR.n505 VGND 0.001416f
C1608 VPWR.n506 VGND 0.005451f
C1609 VPWR.n507 VGND 0.002356f
C1610 VPWR.n508 VGND 0.005451f
C1611 VPWR.t92 VGND 0.002227f
C1612 VPWR.t83 VGND 0.002227f
C1613 VPWR.n509 VGND 0.004781f
C1614 VPWR.n510 VGND 0.001795f
C1615 VPWR.t91 VGND 0.008481f
C1616 VPWR.n511 VGND 0.009967f
C1617 VPWR.n512 VGND 0.004545f
C1618 VPWR.n513 VGND 0.007286f
C1619 VPWR.n514 VGND 0.007286f
C1620 VPWR.n515 VGND 0.001613f
C1621 VPWR.n516 VGND 0.005451f
C1622 VPWR.n517 VGND 0.002258f
C1623 VPWR.n518 VGND 0.001388f
C1624 VPWR.n519 VGND 0.007127f
C1625 VPWR.n520 VGND 0.292827f
C1626 VPWR.n521 VGND 5.29883f
C1627 VPWR.n522 VGND 0.624707f
C1628 VPWR.n523 VGND 0.67635f
C1629 VPWR.n524 VGND 0.110768f
C1630 VPWR.n525 VGND 0.110713f
C1631 VPWR.n526 VGND 0.221562f
C1632 VPWR.n527 VGND 0.221726f
C1633 VPWR.n528 VGND 0.673418f
C1634 VPWR.n529 VGND 0.110658f
C1635 VPWR.n530 VGND 0.111014f
C1636 VPWR.n531 VGND 0.661726f
C1637 VPWR.n532 VGND 0.110363f
C1638 VPWR.n533 VGND 0.110011f
C1639 VPWR.n534 VGND 0.220238f
C1640 VPWR.n535 VGND 0.660872f
C1641 VPWR.n536 VGND 0.675931f
C1642 VPWR.n537 VGND 0.66258f
C1643 VPWR.n538 VGND 0.220458f
C1644 VPWR.n539 VGND 0.110201f
C1645 VPWR.n540 VGND 0.110255f
C1646 VPWR.n541 VGND 0.379109f
C1647 VPWR.n542 VGND 0.707327f
C1648 VPWR.t268 VGND 0.038813f
C1649 VPWR.t270 VGND 0.00879f
C1650 VPWR.n543 VGND 0.05086f
C1651 VPWR.t182 VGND 0.002392f
C1652 VPWR.t168 VGND 0.002392f
C1653 VPWR.n544 VGND 0.004947f
C1654 VPWR.n545 VGND 0.098234f
C1655 VPWR.t170 VGND 0.002392f
C1656 VPWR.t174 VGND 0.002392f
C1657 VPWR.n546 VGND 0.004947f
C1658 VPWR.n547 VGND 0.082582f
C1659 VPWR.t262 VGND 0.038787f
C1660 VPWR.t264 VGND 0.00879f
C1661 VPWR.n548 VGND 0.090806f
C1662 VPWR.t172 VGND 0.002392f
C1663 VPWR.t176 VGND 0.002392f
C1664 VPWR.n549 VGND 0.004947f
C1665 VPWR.n550 VGND 0.119761f
C1666 VPWR.t166 VGND 0.002392f
C1667 VPWR.t184 VGND 0.002392f
C1668 VPWR.n551 VGND 0.004947f
C1669 VPWR.n552 VGND 0.072188f
C1670 VPWR.t269 VGND 0.136425f
C1671 VPWR.t181 VGND 0.108971f
C1672 VPWR.t167 VGND 0.108971f
C1673 VPWR.t169 VGND 0.108971f
C1674 VPWR.t173 VGND 0.108971f
C1675 VPWR.t179 VGND 0.078349f
C1676 VPWR.t263 VGND 0.136425f
C1677 VPWR.t175 VGND 0.108971f
C1678 VPWR.t171 VGND 0.108971f
C1679 VPWR.t183 VGND 0.108971f
C1680 VPWR.t165 VGND 0.108971f
C1681 VPWR.t177 VGND 0.085107f
C1682 VPWR.n553 VGND -0.063904f
C1683 VPWR.t162 VGND 0.091784f
C1684 VPWR.n554 VGND 0.140992f
C1685 VPWR.n555 VGND 0.018809f
C1686 VPWR.t180 VGND 0.002392f
C1687 VPWR.t178 VGND 0.002392f
C1688 VPWR.n556 VGND 0.004947f
C1689 VPWR.n557 VGND 0.081171f
C1690 VPWR.n558 VGND 2.89145f
C1691 VPWR.n559 VGND 1.42069f
C1692 VPWR.n560 VGND 3.70727f
C1693 VPWR.n561 VGND 0.029122f
C1694 VPWR.n562 VGND 0.016784f
C1695 VPWR.n563 VGND 0.119794f
C1696 VPWR.t284 VGND 0.095507f
C1697 VPWR.n564 VGND 0.060445f
C1698 VPWR.t40 VGND 0.095507f
C1699 VPWR.n565 VGND 0.098959f
C1700 VPWR.n566 VGND 0.05179f
C1701 VPWR.n567 VGND 0.228182f
C1702 VPWR.n568 VGND 0.029122f
C1703 VPWR.n569 VGND 0.016784f
C1704 VPWR.n570 VGND 0.119794f
C1705 VPWR.t163 VGND 0.095507f
C1706 VPWR.n571 VGND 0.060445f
C1707 VPWR.t164 VGND 0.095507f
C1708 VPWR.n572 VGND 0.098959f
C1709 VPWR.n573 VGND 0.05179f
C1710 VPWR.n574 VGND 0.23101f
C1711 VPWR.n575 VGND 0.212637f
C1712 VPWR.n576 VGND 2.81733f
C1713 VPWR.n577 VGND 0.003801f
C1714 VPWR.n578 VGND 0.007286f
C1715 VPWR.t45 VGND 0.002227f
C1716 VPWR.t43 VGND 0.002227f
C1717 VPWR.n579 VGND 0.004781f
C1718 VPWR.t42 VGND 0.002227f
C1719 VPWR.t44 VGND 0.002227f
C1720 VPWR.n580 VGND 0.004781f
C1721 VPWR.n581 VGND 0.001991f
C1722 VPWR.t282 VGND 0.00848f
C1723 VPWR.n582 VGND 0.012082f
C1724 VPWR.n583 VGND 0.005464f
C1725 VPWR.n584 VGND 0.007286f
C1726 VPWR.n585 VGND 0.007286f
C1727 VPWR.n586 VGND 0.001416f
C1728 VPWR.n587 VGND 0.005451f
C1729 VPWR.n588 VGND 0.002356f
C1730 VPWR.n589 VGND 0.005451f
C1731 VPWR.t281 VGND 0.002227f
C1732 VPWR.t283 VGND 0.002227f
C1733 VPWR.n590 VGND 0.004781f
C1734 VPWR.n591 VGND 0.001795f
C1735 VPWR.t39 VGND 0.008481f
C1736 VPWR.n592 VGND 0.009967f
C1737 VPWR.n593 VGND 0.004545f
C1738 VPWR.n594 VGND 0.007286f
C1739 VPWR.n595 VGND 0.007286f
C1740 VPWR.n596 VGND 0.001613f
C1741 VPWR.n597 VGND 0.005451f
C1742 VPWR.n598 VGND 0.002258f
C1743 VPWR.n599 VGND 0.001388f
C1744 VPWR.n600 VGND 0.007127f
C1745 VPWR.n601 VGND 0.292827f
C1746 VPWR.n602 VGND 3.83551f
C1747 VPWR.n603 VGND 0.624707f
C1748 VPWR.n604 VGND 0.67635f
C1749 VPWR.n605 VGND 0.110768f
C1750 VPWR.n606 VGND 0.110713f
C1751 VPWR.n607 VGND 0.221562f
C1752 VPWR.n608 VGND 0.221726f
C1753 VPWR.n609 VGND 0.673418f
C1754 VPWR.n610 VGND 0.110658f
C1755 VPWR.n611 VGND 0.111014f
C1756 VPWR.n612 VGND 0.661726f
C1757 VPWR.n613 VGND 0.110363f
C1758 VPWR.n614 VGND 0.110011f
C1759 VPWR.n615 VGND 0.220238f
C1760 VPWR.n616 VGND 0.660872f
C1761 VPWR.n617 VGND 0.675931f
C1762 VPWR.n618 VGND 0.66258f
C1763 VPWR.n619 VGND 0.220458f
C1764 VPWR.n620 VGND 0.110201f
C1765 VPWR.n621 VGND 0.110255f
C1766 VPWR.n622 VGND 0.379109f
C1767 VPWR.n623 VGND 0.707327f
C1768 VPWR.t274 VGND 0.038813f
C1769 VPWR.t276 VGND 0.00879f
C1770 VPWR.n624 VGND 0.05086f
C1771 VPWR.t130 VGND 0.002392f
C1772 VPWR.t120 VGND 0.002392f
C1773 VPWR.n625 VGND 0.004947f
C1774 VPWR.n626 VGND 0.098234f
C1775 VPWR.t118 VGND 0.002392f
C1776 VPWR.t124 VGND 0.002392f
C1777 VPWR.n627 VGND 0.004947f
C1778 VPWR.n628 VGND 0.082582f
C1779 VPWR.t271 VGND 0.038787f
C1780 VPWR.t273 VGND 0.00879f
C1781 VPWR.n629 VGND 0.090806f
C1782 VPWR.t122 VGND 0.002392f
C1783 VPWR.t126 VGND 0.002392f
C1784 VPWR.n630 VGND 0.004947f
C1785 VPWR.n631 VGND 0.119761f
C1786 VPWR.t116 VGND 0.002392f
C1787 VPWR.t114 VGND 0.002392f
C1788 VPWR.n632 VGND 0.004947f
C1789 VPWR.n633 VGND 0.072188f
C1790 VPWR.t275 VGND 0.136425f
C1791 VPWR.t129 VGND 0.108971f
C1792 VPWR.t119 VGND 0.108971f
C1793 VPWR.t117 VGND 0.108971f
C1794 VPWR.t123 VGND 0.108971f
C1795 VPWR.t127 VGND 0.078349f
C1796 VPWR.t272 VGND 0.136425f
C1797 VPWR.t125 VGND 0.108971f
C1798 VPWR.t121 VGND 0.108971f
C1799 VPWR.t113 VGND 0.108971f
C1800 VPWR.t115 VGND 0.108971f
C1801 VPWR.t131 VGND 0.085107f
C1802 VPWR.n634 VGND -0.063904f
C1803 VPWR.t41 VGND 0.091784f
C1804 VPWR.n635 VGND 0.140992f
C1805 VPWR.n636 VGND 0.018809f
C1806 VPWR.t128 VGND 0.002392f
C1807 VPWR.t132 VGND 0.002392f
C1808 VPWR.n637 VGND 0.004947f
C1809 VPWR.n638 VGND 0.081171f
C1810 VPWR.n639 VGND 2.89145f
C1811 VPWR.n640 VGND 1.42069f
C1812 VPWR.n641 VGND 3.70727f
C1813 VPWR.n642 VGND 7.173009f
C1814 ui_in[4].t10 VGND 0.012697f
C1815 ui_in[4].t0 VGND 0.007482f
C1816 ui_in[4].t8 VGND 0.012697f
C1817 ui_in[4].t18 VGND 0.007482f
C1818 ui_in[4].n0 VGND 0.018311f
C1819 ui_in[4].t15 VGND 0.012697f
C1820 ui_in[4].t4 VGND 0.007482f
C1821 ui_in[4].t13 VGND 0.012697f
C1822 ui_in[4].t2 VGND 0.007482f
C1823 ui_in[4].n1 VGND 0.018311f
C1824 ui_in[4].t9 VGND 0.012697f
C1825 ui_in[4].t19 VGND 0.007482f
C1826 ui_in[4].n2 VGND 0.017114f
C1827 ui_in[4].n3 VGND 0.00838f
C1828 ui_in[4].n4 VGND 0.006953f
C1829 ui_in[4].n5 VGND 0.00838f
C1830 ui_in[4].n6 VGND 0.018311f
C1831 ui_in[4].n7 VGND 0.00838f
C1832 ui_in[4].n8 VGND 0.006953f
C1833 ui_in[4].n9 VGND 0.006953f
C1834 ui_in[4].n10 VGND 0.00838f
C1835 ui_in[4].n11 VGND 0.018311f
C1836 ui_in[4].t7 VGND 0.012697f
C1837 ui_in[4].t17 VGND 0.007482f
C1838 ui_in[4].t5 VGND 0.012697f
C1839 ui_in[4].t11 VGND 0.007482f
C1840 ui_in[4].n12 VGND 0.018311f
C1841 ui_in[4].t14 VGND 0.012697f
C1842 ui_in[4].t3 VGND 0.007482f
C1843 ui_in[4].n13 VGND 0.017114f
C1844 ui_in[4].n14 VGND 0.008954f
C1845 ui_in[4].n15 VGND 0.006953f
C1846 ui_in[4].n16 VGND 0.00838f
C1847 ui_in[4].n17 VGND 0.018311f
C1848 ui_in[4].n18 VGND 0.00838f
C1849 ui_in[4].n19 VGND 0.006273f
C1850 ui_in[4].n20 VGND 0.426388f
C1851 ui_in[4].t1 VGND 0.13816f
C1852 ui_in[4].t12 VGND 0.138158f
C1853 ui_in[4].n21 VGND 0.799636f
C1854 ui_in[4].n22 VGND 0.524745f
C1855 ui_in[4].n23 VGND 2.78873f
C1856 ui_in[4].t16 VGND 0.141867f
C1857 ui_in[4].t6 VGND 0.141865f
C1858 ui_in[4].n24 VGND 0.782844f
C1859 ui_in[4].n25 VGND 0.530543f
C1860 ui_in[4].n26 VGND 1.47469f
.ends

