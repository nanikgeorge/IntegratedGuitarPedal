magic
tech sky130A
magscale 1 2
timestamp 1713488381
<< pwell >>
rect -201 -782 201 782
<< psubdiff >>
rect -165 712 -69 746
rect 69 712 165 746
rect -165 650 -131 712
rect 131 650 165 712
rect -165 -712 -131 -650
rect 131 -712 165 -650
rect -165 -746 -69 -712
rect 69 -746 165 -712
<< psubdiffcont >>
rect -69 712 69 746
rect -165 -650 -131 650
rect 131 -650 165 650
rect -69 -746 69 -712
<< xpolycontact >>
rect -35 184 35 616
rect -35 -616 35 -184
<< xpolyres >>
rect -35 -184 35 184
<< locali >>
rect -165 712 -69 746
rect 69 712 165 746
rect -165 650 -131 712
rect 131 650 165 712
rect -165 -712 -131 -650
rect 131 -712 165 -650
rect -165 -746 -69 -712
rect 69 -746 165 -712
<< viali >>
rect -19 201 19 598
rect -19 -598 19 -201
<< metal1 >>
rect -25 598 25 610
rect -25 201 -19 598
rect 19 201 25 598
rect -25 189 25 201
rect -25 -201 25 -189
rect -25 -598 -19 -201
rect 19 -598 25 -201
rect -25 -610 25 -598
<< properties >>
string FIXED_BBOX -148 -729 148 729
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 2 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 12.504k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
