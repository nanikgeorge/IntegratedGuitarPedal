magic
tech sky130A
magscale 1 2
timestamp 1713310215
<< nwell >>
rect 26 512 3252 1024
<< pwell >>
rect 20 -370 3250 -200
<< nmos >>
rect 120 185 320 385
rect 378 185 578 385
rect 636 185 836 385
rect 894 185 1094 385
rect 1152 185 1352 385
rect 1410 185 1610 385
rect 1668 185 1868 385
rect 1926 185 2126 385
rect 2184 185 2384 385
rect 2442 185 2642 385
rect 2700 185 2900 385
rect 2958 185 3158 385
rect 120 -135 320 -51
rect 378 -135 578 -51
rect 636 -135 836 -51
rect 894 -135 1094 -51
rect 1152 -135 1352 -51
rect 1410 -135 1610 -51
rect 1668 -135 1868 -51
rect 1926 -135 2126 -51
rect 2184 -135 2384 -51
rect 2442 -135 2642 -51
rect 2700 -135 2900 -51
rect 2958 -135 3158 -51
<< pmos >>
rect 120 612 320 812
rect 378 612 578 812
rect 636 612 836 812
rect 894 612 1094 812
rect 1152 612 1352 812
rect 1410 612 1610 812
rect 1668 612 1868 812
rect 1926 612 2126 812
rect 2184 612 2384 812
rect 2442 612 2642 812
rect 2700 612 2900 812
rect 2958 612 3158 812
<< ndiff >>
rect 62 373 120 385
rect 62 197 74 373
rect 108 197 120 373
rect 62 185 120 197
rect 320 373 378 385
rect 320 197 332 373
rect 366 197 378 373
rect 320 185 378 197
rect 578 373 636 385
rect 578 197 590 373
rect 624 197 636 373
rect 578 185 636 197
rect 836 373 894 385
rect 836 197 848 373
rect 882 197 894 373
rect 836 185 894 197
rect 1094 373 1152 385
rect 1094 197 1106 373
rect 1140 197 1152 373
rect 1094 185 1152 197
rect 1352 373 1410 385
rect 1352 197 1364 373
rect 1398 197 1410 373
rect 1352 185 1410 197
rect 1610 373 1668 385
rect 1610 197 1622 373
rect 1656 197 1668 373
rect 1610 185 1668 197
rect 1868 373 1926 385
rect 1868 197 1880 373
rect 1914 197 1926 373
rect 1868 185 1926 197
rect 2126 373 2184 385
rect 2126 197 2138 373
rect 2172 197 2184 373
rect 2126 185 2184 197
rect 2384 373 2442 385
rect 2384 197 2396 373
rect 2430 197 2442 373
rect 2384 185 2442 197
rect 2642 373 2700 385
rect 2642 197 2654 373
rect 2688 197 2700 373
rect 2642 185 2700 197
rect 2900 373 2958 385
rect 2900 197 2912 373
rect 2946 197 2958 373
rect 2900 185 2958 197
rect 3158 373 3216 385
rect 3158 197 3170 373
rect 3204 197 3216 373
rect 3158 185 3216 197
rect 62 -63 120 -51
rect 62 -123 74 -63
rect 108 -123 120 -63
rect 62 -135 120 -123
rect 320 -63 378 -51
rect 320 -123 332 -63
rect 366 -123 378 -63
rect 320 -135 378 -123
rect 578 -63 636 -51
rect 578 -123 590 -63
rect 624 -123 636 -63
rect 578 -135 636 -123
rect 836 -63 894 -51
rect 836 -123 848 -63
rect 882 -123 894 -63
rect 836 -135 894 -123
rect 1094 -63 1152 -51
rect 1094 -123 1106 -63
rect 1140 -123 1152 -63
rect 1094 -135 1152 -123
rect 1352 -63 1410 -51
rect 1352 -123 1364 -63
rect 1398 -123 1410 -63
rect 1352 -135 1410 -123
rect 1610 -63 1668 -51
rect 1610 -123 1622 -63
rect 1656 -123 1668 -63
rect 1610 -135 1668 -123
rect 1868 -63 1926 -51
rect 1868 -123 1880 -63
rect 1914 -123 1926 -63
rect 1868 -135 1926 -123
rect 2126 -63 2184 -51
rect 2126 -123 2138 -63
rect 2172 -123 2184 -63
rect 2126 -135 2184 -123
rect 2384 -63 2442 -51
rect 2384 -123 2396 -63
rect 2430 -123 2442 -63
rect 2384 -135 2442 -123
rect 2642 -63 2700 -51
rect 2642 -123 2654 -63
rect 2688 -123 2700 -63
rect 2642 -135 2700 -123
rect 2900 -63 2958 -51
rect 2900 -123 2912 -63
rect 2946 -123 2958 -63
rect 2900 -135 2958 -123
rect 3158 -63 3216 -51
rect 3158 -123 3170 -63
rect 3204 -123 3216 -63
rect 3158 -135 3216 -123
<< pdiff >>
rect 62 800 120 812
rect 62 624 74 800
rect 108 624 120 800
rect 62 612 120 624
rect 320 800 378 812
rect 320 624 332 800
rect 366 624 378 800
rect 320 612 378 624
rect 578 800 636 812
rect 578 624 590 800
rect 624 624 636 800
rect 578 612 636 624
rect 836 800 894 812
rect 836 624 848 800
rect 882 624 894 800
rect 836 612 894 624
rect 1094 800 1152 812
rect 1094 624 1106 800
rect 1140 624 1152 800
rect 1094 612 1152 624
rect 1352 800 1410 812
rect 1352 624 1364 800
rect 1398 624 1410 800
rect 1352 612 1410 624
rect 1610 800 1668 812
rect 1610 624 1622 800
rect 1656 624 1668 800
rect 1610 612 1668 624
rect 1868 800 1926 812
rect 1868 624 1880 800
rect 1914 624 1926 800
rect 1868 612 1926 624
rect 2126 800 2184 812
rect 2126 624 2138 800
rect 2172 624 2184 800
rect 2126 612 2184 624
rect 2384 800 2442 812
rect 2384 624 2396 800
rect 2430 624 2442 800
rect 2384 612 2442 624
rect 2642 800 2700 812
rect 2642 624 2654 800
rect 2688 624 2700 800
rect 2642 612 2700 624
rect 2900 800 2958 812
rect 2900 624 2912 800
rect 2946 624 2958 800
rect 2900 612 2958 624
rect 3158 800 3216 812
rect 3158 624 3170 800
rect 3204 624 3216 800
rect 3158 612 3216 624
<< ndiffc >>
rect 74 197 108 373
rect 332 197 366 373
rect 590 197 624 373
rect 848 197 882 373
rect 1106 197 1140 373
rect 1364 197 1398 373
rect 1622 197 1656 373
rect 1880 197 1914 373
rect 2138 197 2172 373
rect 2396 197 2430 373
rect 2654 197 2688 373
rect 2912 197 2946 373
rect 3170 197 3204 373
rect 74 -123 108 -63
rect 332 -123 366 -63
rect 590 -123 624 -63
rect 848 -123 882 -63
rect 1106 -123 1140 -63
rect 1364 -123 1398 -63
rect 1622 -123 1656 -63
rect 1880 -123 1914 -63
rect 2138 -123 2172 -63
rect 2396 -123 2430 -63
rect 2654 -123 2688 -63
rect 2912 -123 2946 -63
rect 3170 -123 3204 -63
<< pdiffc >>
rect 74 624 108 800
rect 332 624 366 800
rect 590 624 624 800
rect 848 624 882 800
rect 1106 624 1140 800
rect 1364 624 1398 800
rect 1622 624 1656 800
rect 1880 624 1914 800
rect 2138 624 2172 800
rect 2396 624 2430 800
rect 2654 624 2688 800
rect 2912 624 2946 800
rect 3170 624 3204 800
<< psubdiff >>
rect 70 -250 3200 -220
rect 70 -300 110 -250
rect 3160 -300 3200 -250
rect 70 -329 3200 -300
rect 70 -330 430 -329
rect 2840 -330 3200 -329
<< nsubdiff >>
rect 110 940 3200 980
rect 110 900 150 940
rect 3160 900 3200 940
rect 110 870 3200 900
<< psubdiffcont >>
rect 110 -300 3160 -250
<< nsubdiffcont >>
rect 150 900 3160 940
<< poly >>
rect 120 812 320 838
rect 378 812 578 838
rect 636 812 836 838
rect 894 812 1094 838
rect 1152 812 1352 838
rect 1410 812 1610 838
rect 1668 812 1868 838
rect 1926 812 2126 838
rect 2184 812 2384 838
rect 2442 812 2642 838
rect 2700 812 2900 838
rect 2958 812 3158 838
rect 120 565 320 612
rect 120 531 136 565
rect 304 531 320 565
rect 120 515 320 531
rect 378 565 578 612
rect 378 531 394 565
rect 562 531 578 565
rect 378 515 578 531
rect 636 565 836 612
rect 636 531 652 565
rect 820 531 836 565
rect 636 515 836 531
rect 894 565 1094 612
rect 894 531 910 565
rect 1078 531 1094 565
rect 894 515 1094 531
rect 1152 565 1352 612
rect 1152 531 1168 565
rect 1336 531 1352 565
rect 1152 515 1352 531
rect 1410 565 1610 612
rect 1410 531 1426 565
rect 1594 531 1610 565
rect 1410 515 1610 531
rect 1668 565 1868 612
rect 1668 531 1684 565
rect 1852 531 1868 565
rect 1668 515 1868 531
rect 1926 565 2126 612
rect 1926 531 1942 565
rect 2110 531 2126 565
rect 1926 515 2126 531
rect 2184 565 2384 612
rect 2184 531 2200 565
rect 2368 531 2384 565
rect 2184 515 2384 531
rect 2442 565 2642 612
rect 2442 531 2458 565
rect 2626 531 2642 565
rect 2442 515 2642 531
rect 2700 565 2900 612
rect 2700 531 2716 565
rect 2884 531 2900 565
rect 2700 515 2900 531
rect 2958 565 3158 612
rect 2958 531 2974 565
rect 3142 531 3158 565
rect 2958 515 3158 531
rect 378 457 578 473
rect 378 423 394 457
rect 562 423 578 457
rect 120 385 320 411
rect 378 385 578 423
rect 1152 457 1352 473
rect 1152 423 1168 457
rect 1336 423 1352 457
rect 636 385 836 411
rect 894 385 1094 411
rect 1152 385 1352 423
rect 1410 457 1610 473
rect 1410 423 1426 457
rect 1594 423 1610 457
rect 1410 385 1610 423
rect 2184 457 2384 473
rect 2184 423 2200 457
rect 2368 423 2384 457
rect 1668 385 1868 411
rect 1926 385 2126 411
rect 2184 385 2384 423
rect 2442 457 2642 473
rect 2442 423 2458 457
rect 2626 423 2642 457
rect 2442 385 2642 423
rect 2700 385 2900 411
rect 2958 385 3158 411
rect 120 147 320 185
rect 378 159 578 185
rect 120 113 136 147
rect 304 113 320 147
rect 120 97 320 113
rect 636 147 836 185
rect 636 113 652 147
rect 820 113 836 147
rect 636 97 836 113
rect 894 147 1094 185
rect 1152 159 1352 185
rect 1410 159 1610 185
rect 894 113 910 147
rect 1078 113 1094 147
rect 894 97 1094 113
rect 1668 147 1868 185
rect 1668 113 1684 147
rect 1852 113 1868 147
rect 1668 97 1868 113
rect 1926 147 2126 185
rect 2184 159 2384 185
rect 2442 159 2642 185
rect 1926 113 1942 147
rect 2110 113 2126 147
rect 1926 97 2126 113
rect 2700 147 2900 185
rect 2700 113 2716 147
rect 2884 113 2900 147
rect 2700 97 2900 113
rect 2958 147 3158 185
rect 2958 113 2974 147
rect 3142 113 3158 147
rect 2958 97 3158 113
rect 120 21 320 37
rect 120 -13 136 21
rect 304 -13 320 21
rect 120 -51 320 -13
rect 378 21 578 37
rect 378 -13 394 21
rect 562 -13 578 21
rect 378 -51 578 -13
rect 636 21 836 37
rect 636 -13 652 21
rect 820 -13 836 21
rect 636 -51 836 -13
rect 894 21 1094 37
rect 894 -13 910 21
rect 1078 -13 1094 21
rect 894 -51 1094 -13
rect 1152 21 1352 37
rect 1152 -13 1168 21
rect 1336 -13 1352 21
rect 1152 -51 1352 -13
rect 1410 21 1610 37
rect 1410 -13 1426 21
rect 1594 -13 1610 21
rect 1410 -51 1610 -13
rect 1668 21 1868 37
rect 1668 -13 1684 21
rect 1852 -13 1868 21
rect 1668 -51 1868 -13
rect 1926 21 2126 37
rect 1926 -13 1942 21
rect 2110 -13 2126 21
rect 1926 -51 2126 -13
rect 2184 21 2384 37
rect 2184 -13 2200 21
rect 2368 -13 2384 21
rect 2184 -51 2384 -13
rect 2442 21 2642 37
rect 2442 -13 2458 21
rect 2626 -13 2642 21
rect 2442 -51 2642 -13
rect 2700 21 2900 37
rect 2700 -13 2716 21
rect 2884 -13 2900 21
rect 2700 -51 2900 -13
rect 2958 21 3158 37
rect 2958 -13 2974 21
rect 3142 -13 3158 21
rect 2958 -51 3158 -13
rect 120 -161 320 -135
rect 378 -161 578 -135
rect 636 -161 836 -135
rect 894 -161 1094 -135
rect 1152 -161 1352 -135
rect 1410 -161 1610 -135
rect 1668 -161 1868 -135
rect 1926 -161 2126 -135
rect 2184 -161 2384 -135
rect 2442 -161 2642 -135
rect 2700 -161 2900 -135
rect 2958 -161 3158 -135
<< polycont >>
rect 136 531 304 565
rect 394 531 562 565
rect 652 531 820 565
rect 910 531 1078 565
rect 1168 531 1336 565
rect 1426 531 1594 565
rect 1684 531 1852 565
rect 1942 531 2110 565
rect 2200 531 2368 565
rect 2458 531 2626 565
rect 2716 531 2884 565
rect 2974 531 3142 565
rect 394 423 562 457
rect 1168 423 1336 457
rect 1426 423 1594 457
rect 2200 423 2368 457
rect 2458 423 2626 457
rect 136 113 304 147
rect 652 113 820 147
rect 910 113 1078 147
rect 1684 113 1852 147
rect 1942 113 2110 147
rect 2716 113 2884 147
rect 2974 113 3142 147
rect 136 -13 304 21
rect 394 -13 562 21
rect 652 -13 820 21
rect 910 -13 1078 21
rect 1168 -13 1336 21
rect 1426 -13 1594 21
rect 1684 -13 1852 21
rect 1942 -13 2110 21
rect 2200 -13 2368 21
rect 2458 -13 2626 21
rect 2716 -13 2884 21
rect 2974 -13 3142 21
<< locali >>
rect -480 940 3210 980
rect -480 900 -420 940
rect 3160 900 3210 940
rect -480 860 3210 900
rect 74 800 108 816
rect 74 608 108 624
rect 332 800 366 816
rect 332 608 366 624
rect 590 800 624 816
rect 590 608 624 624
rect 848 800 882 816
rect 848 608 882 624
rect 1106 800 1140 816
rect 1106 608 1140 624
rect 1364 800 1398 816
rect 1364 608 1398 624
rect 1622 800 1656 816
rect 1622 608 1656 624
rect 1880 800 1914 816
rect 1880 608 1914 624
rect 2138 800 2172 816
rect 2138 608 2172 624
rect 2396 800 2430 816
rect 2396 608 2430 624
rect 2654 800 2688 816
rect 2654 608 2688 624
rect 2912 800 2946 816
rect 2912 608 2946 624
rect 3170 800 3204 816
rect 3170 608 3204 624
rect 120 531 136 565
rect 304 531 320 565
rect 378 531 394 565
rect 562 531 578 565
rect 636 531 652 565
rect 820 531 836 565
rect 894 531 910 565
rect 1078 531 1094 565
rect 1152 531 1168 565
rect 1336 531 1352 565
rect 1410 531 1426 565
rect 1594 531 1610 565
rect 1668 531 1684 565
rect 1852 531 1868 565
rect 1926 531 1942 565
rect 2110 531 2126 565
rect 2184 531 2200 565
rect 2368 531 2384 565
rect 2442 531 2458 565
rect 2626 531 2642 565
rect 2700 531 2716 565
rect 2884 531 2900 565
rect 2958 531 2974 565
rect 3142 531 3158 565
rect 378 423 394 457
rect 562 423 578 457
rect 1152 423 1168 457
rect 1336 423 1352 457
rect 1410 423 1426 457
rect 1594 423 1610 457
rect 2184 423 2200 457
rect 2368 423 2384 457
rect 2442 423 2458 457
rect 2626 423 2642 457
rect 74 373 108 389
rect 74 181 108 197
rect 332 373 366 389
rect 332 181 366 197
rect 590 373 624 389
rect 590 181 624 197
rect 848 373 882 389
rect 848 181 882 197
rect 1106 373 1140 389
rect 1106 181 1140 197
rect 1364 373 1398 389
rect 1364 181 1398 197
rect 1622 373 1656 389
rect 1622 181 1656 197
rect 1880 373 1914 389
rect 1880 181 1914 197
rect 2138 373 2172 389
rect 2138 181 2172 197
rect 2396 373 2430 389
rect 2396 181 2430 197
rect 2654 373 2688 389
rect 2654 181 2688 197
rect 2912 373 2946 389
rect 2912 181 2946 197
rect 3170 373 3204 389
rect 3170 181 3204 197
rect 120 113 136 147
rect 304 113 320 147
rect 636 113 652 147
rect 820 113 836 147
rect 894 113 910 147
rect 1078 113 1094 147
rect 1668 113 1684 147
rect 1852 113 1868 147
rect 1926 113 1942 147
rect 2110 113 2126 147
rect 2700 113 2716 147
rect 2884 113 2900 147
rect 2958 113 2974 147
rect 3142 113 3158 147
rect 120 -13 136 21
rect 304 -13 320 21
rect 378 -13 394 21
rect 562 -13 578 21
rect 636 -13 652 21
rect 820 -13 836 21
rect 894 -13 910 21
rect 1078 -13 1094 21
rect 1152 -13 1168 21
rect 1336 -13 1352 21
rect 1410 -13 1426 21
rect 1594 -13 1610 21
rect 1668 -13 1684 21
rect 1852 -13 1868 21
rect 1926 -13 1942 21
rect 2110 -13 2126 21
rect 2184 -13 2200 21
rect 2368 -13 2384 21
rect 2442 -13 2458 21
rect 2626 -13 2642 21
rect 2700 -13 2716 21
rect 2884 -13 2900 21
rect 2958 -13 2974 21
rect 3142 -13 3158 21
rect 74 -63 108 -47
rect 74 -139 108 -123
rect 332 -63 366 -47
rect 332 -139 366 -123
rect 590 -63 624 -47
rect 590 -139 624 -123
rect 848 -63 882 -47
rect 848 -139 882 -123
rect 1106 -63 1140 -47
rect 1106 -139 1140 -123
rect 1364 -63 1398 -47
rect 1364 -139 1398 -123
rect 1622 -63 1656 -47
rect 1622 -139 1656 -123
rect 1880 -63 1914 -47
rect 1880 -139 1914 -123
rect 2138 -63 2172 -47
rect 2138 -139 2172 -123
rect 2396 -63 2430 -47
rect 2396 -139 2430 -123
rect 2654 -63 2688 -47
rect 2654 -139 2688 -123
rect 2912 -63 2946 -47
rect 2912 -139 2946 -123
rect 3170 -63 3204 -47
rect 3170 -139 3204 -123
rect -480 -190 -40 -160
rect -480 -280 -460 -190
rect -60 -280 -40 -190
rect -480 -300 -40 -280
rect 70 -250 3210 -220
rect 70 -300 110 -250
rect 3160 -300 3210 -250
rect 70 -330 3210 -300
<< viali >>
rect -420 900 150 940
rect 150 900 3160 940
rect 74 624 108 800
rect 332 624 366 800
rect 590 624 624 800
rect 848 624 882 800
rect 1106 624 1140 800
rect 1364 624 1398 800
rect 1622 624 1656 800
rect 1880 624 1914 800
rect 2138 624 2172 800
rect 2396 624 2430 800
rect 2654 624 2688 800
rect 2912 624 2946 800
rect 3170 624 3204 800
rect 136 531 304 565
rect 394 531 562 565
rect 652 531 820 565
rect 910 531 1078 565
rect 1168 531 1336 565
rect 1426 531 1594 565
rect 1684 531 1852 565
rect 1942 531 2110 565
rect 2200 531 2368 565
rect 2458 531 2626 565
rect 2716 531 2884 565
rect 2974 531 3142 565
rect 394 423 562 457
rect 1168 423 1336 457
rect 1426 423 1594 457
rect 2200 423 2368 457
rect 2458 423 2626 457
rect 74 197 108 373
rect 332 197 366 373
rect 590 197 624 373
rect 848 197 882 373
rect 1106 197 1140 373
rect 1364 197 1398 373
rect 1622 197 1656 373
rect 1880 197 1914 373
rect 2138 197 2172 373
rect 2396 197 2430 373
rect 2654 197 2688 373
rect 2912 197 2946 373
rect 3170 197 3204 373
rect 136 113 304 147
rect 652 113 820 147
rect 910 113 1078 147
rect 1684 113 1852 147
rect 1942 113 2110 147
rect 2716 113 2884 147
rect 2974 113 3142 147
rect 136 -13 304 21
rect 394 -13 562 21
rect 652 -13 820 21
rect 910 -13 1078 21
rect 1168 -13 1336 21
rect 1426 -13 1594 21
rect 1684 -13 1852 21
rect 1942 -13 2110 21
rect 2200 -13 2368 21
rect 2458 -13 2626 21
rect 2716 -13 2884 21
rect 2974 -13 3142 21
rect 74 -123 108 -63
rect 332 -123 366 -63
rect 590 -123 624 -63
rect 848 -123 882 -63
rect 1106 -123 1140 -63
rect 1364 -123 1398 -63
rect 1622 -123 1656 -63
rect 1880 -123 1914 -63
rect 2138 -123 2172 -63
rect 2396 -123 2430 -63
rect 2654 -123 2688 -63
rect 2912 -123 2946 -63
rect 3170 -123 3204 -63
rect -460 -280 -60 -190
rect 110 -300 3160 -250
<< metal1 >>
rect -480 960 3210 980
rect -480 940 30 960
rect -480 900 -420 940
rect -480 880 30 900
rect 3190 880 3210 960
rect -480 860 3210 880
rect 70 812 130 860
rect 68 800 130 812
rect 320 810 380 820
rect 68 624 74 800
rect 108 624 130 800
rect 68 612 130 624
rect 280 800 430 810
rect 280 690 332 800
rect 366 690 430 800
rect 280 630 290 690
rect 400 630 430 690
rect 280 624 332 630
rect 366 624 430 630
rect 280 620 430 624
rect 540 800 670 860
rect 842 810 888 812
rect 540 624 590 800
rect 624 624 670 800
rect 540 620 670 624
rect 800 800 930 810
rect 800 690 848 800
rect 882 690 930 800
rect 800 630 810 690
rect 920 630 930 690
rect 800 624 848 630
rect 882 624 930 630
rect 800 620 930 624
rect 1060 800 1190 860
rect 1060 624 1106 800
rect 1140 624 1190 800
rect 1060 620 1190 624
rect 1310 800 1440 820
rect 1310 690 1364 800
rect 1398 690 1440 800
rect 70 571 130 612
rect 320 610 430 620
rect 584 612 630 620
rect 842 612 888 620
rect 1100 612 1146 620
rect 380 571 430 610
rect 1310 580 1320 690
rect 1430 580 1440 690
rect 1570 800 1700 860
rect 1874 810 1920 812
rect 1570 624 1622 800
rect 1656 624 1700 800
rect 1570 620 1700 624
rect 1830 800 1960 810
rect 1830 700 1880 800
rect 1914 700 1960 800
rect 1830 630 1840 700
rect 1950 630 1960 700
rect 1830 624 1880 630
rect 1914 624 1960 630
rect 1830 620 1960 624
rect 2090 800 2220 860
rect 2090 624 2138 800
rect 2172 624 2220 800
rect 2090 620 2220 624
rect 2350 800 2480 820
rect 2350 700 2396 800
rect 2430 700 2480 800
rect 1616 612 1662 620
rect 1874 612 1920 620
rect 2132 612 2178 620
rect 1310 571 1440 580
rect 2350 580 2360 700
rect 2470 580 2480 700
rect 2610 800 2740 860
rect 3170 812 3210 860
rect 2906 810 2952 812
rect 2610 624 2654 800
rect 2688 624 2740 800
rect 2610 620 2740 624
rect 2860 800 2990 810
rect 2860 700 2912 800
rect 2946 700 2990 800
rect 2860 630 2870 700
rect 2980 630 2990 700
rect 2860 624 2912 630
rect 2946 624 2990 630
rect 2860 620 2990 624
rect 3164 800 3210 812
rect 3164 624 3170 800
rect 3204 624 3210 800
rect 2648 612 2694 620
rect 2906 612 2952 620
rect 3164 612 3210 624
rect 3170 580 3210 612
rect 2350 571 2480 580
rect 70 570 316 571
rect 70 565 320 570
rect 380 565 574 571
rect 640 565 832 571
rect 898 565 1090 571
rect 1156 565 1606 571
rect 1672 565 1864 571
rect 1930 565 2122 571
rect 2188 565 2638 571
rect 2704 565 2896 571
rect 2960 565 3210 580
rect 70 531 136 565
rect 304 531 320 565
rect 378 531 394 565
rect 562 531 652 565
rect 820 531 910 565
rect 1078 531 1168 565
rect 1336 531 1426 565
rect 1594 531 1684 565
rect 1852 531 1942 565
rect 2110 531 2200 565
rect 2368 531 2458 565
rect 2626 531 2716 565
rect 2884 531 2900 565
rect 2960 531 2974 565
rect 3142 531 3210 565
rect 70 530 320 531
rect 380 530 574 531
rect 124 525 316 530
rect 382 525 574 530
rect 640 525 832 531
rect 898 525 1090 531
rect 1156 525 1348 531
rect 1414 525 1606 531
rect 1672 525 1864 531
rect 1930 525 2122 531
rect 2188 525 2380 531
rect 2446 525 2638 531
rect 2704 525 2896 531
rect 2960 530 3210 531
rect 2962 525 3154 530
rect 660 480 770 490
rect 382 457 574 463
rect 660 457 670 480
rect 378 423 394 457
rect 562 423 670 457
rect 382 417 574 423
rect 70 385 120 390
rect 68 373 120 385
rect 326 380 372 385
rect 68 197 74 373
rect 108 197 120 373
rect 68 185 120 197
rect 280 373 410 380
rect 280 370 332 373
rect 366 370 410 373
rect 280 310 290 370
rect 400 310 410 370
rect 280 197 332 310
rect 366 197 410 310
rect 584 373 630 385
rect 584 280 590 373
rect 280 190 410 197
rect 540 260 590 280
rect 624 280 630 373
rect 660 320 670 423
rect 760 457 770 480
rect 2730 480 2830 490
rect 1156 457 1348 463
rect 1414 457 1606 463
rect 2188 457 2380 463
rect 2446 457 2638 463
rect 760 423 1168 457
rect 1336 423 1426 457
rect 1594 423 2200 457
rect 2368 423 2458 457
rect 2626 423 2642 457
rect 760 320 770 423
rect 1156 417 1348 423
rect 1414 417 1606 423
rect 2188 417 2380 423
rect 2446 417 2638 423
rect 842 380 888 385
rect 1100 380 1146 385
rect 1358 380 1404 385
rect 1616 380 1662 385
rect 1874 380 1920 385
rect 2132 380 2178 385
rect 2390 380 2436 385
rect 660 310 770 320
rect 800 373 930 380
rect 800 370 848 373
rect 882 370 930 373
rect 800 310 810 370
rect 920 310 930 370
rect 624 260 670 280
rect 540 200 550 260
rect 660 200 670 260
rect 540 197 590 200
rect 624 197 670 200
rect 540 190 670 197
rect 800 197 848 310
rect 882 197 930 310
rect 800 190 930 197
rect 1060 373 1190 380
rect 1060 260 1106 373
rect 1140 260 1190 373
rect 1060 200 1070 260
rect 1180 200 1190 260
rect 1060 197 1106 200
rect 1140 197 1190 200
rect 1060 190 1190 197
rect 1310 373 1440 380
rect 1310 370 1364 373
rect 1398 370 1440 373
rect 1310 310 1320 370
rect 1430 310 1440 370
rect 1310 197 1364 310
rect 1398 197 1440 310
rect 1310 190 1440 197
rect 1580 373 1710 380
rect 1580 260 1622 373
rect 1656 260 1710 373
rect 1580 200 1590 260
rect 1700 200 1710 260
rect 1580 197 1622 200
rect 1656 197 1710 200
rect 1580 190 1710 197
rect 1830 373 1960 380
rect 1830 370 1880 373
rect 1914 370 1960 373
rect 1830 310 1840 370
rect 1950 310 1960 370
rect 1830 197 1880 310
rect 1914 197 1960 310
rect 1830 190 1960 197
rect 2090 373 2220 380
rect 2090 260 2138 373
rect 2172 260 2220 373
rect 2090 200 2100 260
rect 2210 200 2220 260
rect 2090 197 2138 200
rect 2172 197 2220 200
rect 2090 190 2220 197
rect 2350 373 2480 380
rect 2350 370 2396 373
rect 2430 370 2480 373
rect 2350 310 2360 370
rect 2470 310 2480 370
rect 2350 197 2396 310
rect 2430 197 2480 310
rect 2648 373 2694 385
rect 2648 270 2654 373
rect 2350 190 2480 197
rect 2600 260 2654 270
rect 2688 270 2694 373
rect 2730 330 2740 480
rect 2820 330 2830 480
rect 2906 380 2952 385
rect 2730 300 2830 330
rect 2688 260 2730 270
rect 2600 200 2610 260
rect 2720 200 2730 260
rect 2600 197 2654 200
rect 2688 197 2730 200
rect 2600 190 2730 197
rect 326 185 372 190
rect 584 185 630 190
rect 842 185 888 190
rect 1100 185 1146 190
rect 1358 185 1404 190
rect 1616 185 1662 190
rect 1874 185 1920 190
rect 2132 185 2178 190
rect 2390 185 2436 190
rect 2648 185 2694 190
rect 70 180 120 185
rect 70 153 140 180
rect 2760 153 2830 300
rect 2860 373 2990 380
rect 2860 370 2912 373
rect 2946 370 2990 373
rect 2860 310 2870 370
rect 2980 310 2990 370
rect 2860 197 2912 310
rect 2946 197 2990 310
rect 2860 190 2990 197
rect 3160 373 3210 390
rect 3160 197 3170 373
rect 3204 197 3210 373
rect 2906 185 2952 190
rect 3160 180 3210 197
rect 3130 153 3210 180
rect 70 150 316 153
rect 70 147 320 150
rect 640 147 832 153
rect 898 147 1090 153
rect 1672 147 1864 153
rect 1930 147 2122 153
rect 2704 147 2896 153
rect 2962 150 3210 153
rect 2950 147 3210 150
rect 70 113 136 147
rect 304 113 320 147
rect 636 113 652 147
rect 820 113 910 147
rect 1078 113 1684 147
rect 1852 113 1942 147
rect 2110 113 2716 147
rect 2884 113 2900 147
rect 2950 113 2974 147
rect 3142 113 3210 147
rect 70 50 320 113
rect 640 107 832 113
rect 898 107 1090 113
rect 1672 107 1864 113
rect 1930 107 2122 113
rect 2704 107 2896 113
rect 70 21 840 50
rect 1520 40 1530 70
rect 70 -13 136 21
rect 304 -13 394 21
rect 562 -13 652 21
rect 820 -13 840 21
rect 70 -47 840 -13
rect 890 21 1530 40
rect 1750 40 1760 70
rect 2950 50 3210 113
rect 1750 21 2390 40
rect 890 -13 910 21
rect 1078 -13 1168 21
rect 1336 -13 1426 21
rect 1594 -13 1684 10
rect 1852 -13 1942 21
rect 2110 -13 2200 21
rect 2368 -13 2390 21
rect 890 -19 2390 -13
rect 2440 21 3210 50
rect 2440 -13 2458 21
rect 2626 -13 2716 21
rect 2884 -13 2974 21
rect 3142 -13 3210 21
rect 1520 -30 1760 -19
rect 70 -51 884 -47
rect 68 -63 888 -51
rect 68 -123 74 -63
rect 108 -123 332 -63
rect 366 -123 590 -63
rect 624 -123 848 -63
rect 882 -123 888 -63
rect 68 -135 888 -123
rect 1080 -125 1095 -47
rect 1150 -125 1170 -47
rect 1080 -135 1170 -125
rect 1310 -63 1450 -48
rect 1310 -123 1364 -63
rect 1398 -123 1450 -63
rect -480 -170 -40 -160
rect -480 -290 -470 -170
rect -50 -290 -40 -170
rect -480 -300 -40 -290
rect 70 -220 884 -135
rect 1310 -220 1450 -123
rect 1595 -63 1685 -30
rect 1595 -123 1622 -63
rect 1656 -123 1685 -63
rect 1595 -140 1685 -123
rect 1830 -63 1970 -48
rect 1830 -123 1880 -63
rect 1914 -123 1970 -63
rect 1830 -220 1970 -123
rect 2115 -125 2125 -48
rect 2180 -125 2190 -48
rect 2440 -50 3210 -13
rect 2115 -135 2190 -125
rect 2390 -63 3210 -50
rect 2390 -123 2396 -63
rect 2430 -123 2654 -63
rect 2688 -123 2912 -63
rect 2946 -123 3170 -63
rect 3204 -123 3210 -63
rect 2390 -220 3210 -123
rect 70 -240 3210 -220
rect 70 -310 90 -240
rect 3190 -310 3210 -240
rect 70 -330 3210 -310
<< via1 >>
rect 30 940 3190 960
rect 30 900 3160 940
rect 3160 900 3190 940
rect 30 880 3190 900
rect 290 630 332 690
rect 332 630 366 690
rect 366 630 400 690
rect 810 630 848 690
rect 848 630 882 690
rect 882 630 920 690
rect 1320 624 1364 690
rect 1364 624 1398 690
rect 1398 624 1430 690
rect 1320 580 1430 624
rect 1840 630 1880 700
rect 1880 630 1914 700
rect 1914 630 1950 700
rect 2360 624 2396 700
rect 2396 624 2430 700
rect 2430 624 2470 700
rect 2360 580 2470 624
rect 2870 630 2912 700
rect 2912 630 2946 700
rect 2946 630 2980 700
rect 290 310 332 370
rect 332 310 366 370
rect 366 310 400 370
rect 670 320 760 480
rect 810 310 848 370
rect 848 310 882 370
rect 882 310 920 370
rect 550 200 590 260
rect 590 200 624 260
rect 624 200 660 260
rect 1070 200 1106 260
rect 1106 200 1140 260
rect 1140 200 1180 260
rect 1320 310 1364 370
rect 1364 310 1398 370
rect 1398 310 1430 370
rect 1590 200 1622 260
rect 1622 200 1656 260
rect 1656 200 1700 260
rect 1840 310 1880 370
rect 1880 310 1914 370
rect 1914 310 1950 370
rect 2100 200 2138 260
rect 2138 200 2172 260
rect 2172 200 2210 260
rect 2360 310 2396 370
rect 2396 310 2430 370
rect 2430 310 2470 370
rect 2740 330 2820 480
rect 2610 200 2654 260
rect 2654 200 2688 260
rect 2688 200 2720 260
rect 2870 310 2912 370
rect 2912 310 2946 370
rect 2946 310 2980 370
rect 1530 21 1750 70
rect 1530 10 1594 21
rect 1594 10 1684 21
rect 1684 10 1750 21
rect 1095 -63 1150 -47
rect 1095 -123 1106 -63
rect 1106 -123 1140 -63
rect 1140 -123 1150 -63
rect 1095 -125 1150 -123
rect -470 -190 -50 -170
rect -470 -280 -460 -190
rect -460 -280 -60 -190
rect -60 -280 -50 -190
rect -470 -290 -50 -280
rect 2125 -63 2180 -48
rect 2125 -123 2138 -63
rect 2138 -123 2172 -63
rect 2172 -123 2180 -63
rect 2125 -125 2180 -123
rect 90 -250 3190 -240
rect 90 -300 110 -250
rect 110 -300 3160 -250
rect 3160 -300 3190 -250
rect 90 -310 3190 -300
<< metal2 >>
rect 10 1120 3260 1164
rect 10 850 20 1120
rect 3250 850 3260 1120
rect 10 840 3260 850
rect 280 690 410 700
rect 280 630 290 690
rect 400 630 410 690
rect 280 380 410 630
rect 280 310 290 380
rect 400 310 410 380
rect 280 300 410 310
rect 440 690 770 700
rect 440 470 450 690
rect 720 480 770 690
rect 440 320 670 470
rect 760 320 770 480
rect 440 300 770 320
rect 800 690 930 700
rect 800 620 810 690
rect 920 620 930 690
rect 800 370 930 620
rect 800 310 810 370
rect 920 310 930 370
rect 800 300 930 310
rect 1310 690 1440 710
rect 1310 580 1320 690
rect 1430 580 1440 690
rect 1310 380 1440 580
rect 1310 310 1320 380
rect 1430 310 1440 380
rect 1310 300 1440 310
rect 1830 700 1960 710
rect 1830 620 1840 700
rect 1950 620 1960 700
rect 1830 370 1960 620
rect 1830 310 1840 370
rect 1950 310 1960 370
rect 1830 300 1960 310
rect 2350 700 2480 710
rect 2350 580 2360 700
rect 2470 580 2480 700
rect 2350 380 2480 580
rect 2860 700 2990 710
rect 2860 620 2870 700
rect 2980 620 2990 700
rect 2350 310 2360 380
rect 2470 310 2480 380
rect 2530 490 2830 500
rect 2530 320 2550 490
rect 2820 320 2830 490
rect 2530 310 2830 320
rect 2860 370 2990 620
rect 2860 310 2870 370
rect 2980 310 2990 370
rect 2350 300 2480 310
rect 2860 300 2990 310
rect 530 260 2740 270
rect 530 200 550 260
rect 660 200 1070 260
rect 1180 200 1590 260
rect 1700 200 2100 260
rect 2210 200 2610 260
rect 2720 200 2740 260
rect 530 180 2740 200
rect -480 70 1780 110
rect -480 10 1530 70
rect 1750 10 1780 70
rect -480 0 1780 10
rect -480 -170 -40 0
rect 1850 -35 2210 180
rect 1060 -47 2210 -35
rect 1060 -125 1095 -47
rect 1150 -48 2210 -47
rect 1150 -125 2125 -48
rect 2180 -125 2210 -48
rect 1060 -140 2210 -125
rect -480 -290 -470 -170
rect -50 -290 -40 -170
rect -480 -300 -40 -290
rect 10 -450 30 -200
rect 3240 -450 3260 -200
rect 10 -568 3260 -450
<< via2 >>
rect 20 960 3250 1120
rect 20 880 30 960
rect 30 880 3190 960
rect 3190 880 3250 960
rect 20 850 3250 880
rect 290 370 400 380
rect 290 310 400 370
rect 450 480 720 690
rect 450 470 670 480
rect 670 470 720 480
rect 810 630 920 690
rect 810 620 920 630
rect 1320 370 1430 380
rect 1320 310 1430 370
rect 1840 630 1950 690
rect 1840 620 1950 630
rect 2870 630 2980 690
rect 2870 620 2980 630
rect 2360 370 2470 380
rect 2360 310 2470 370
rect 2550 480 2820 490
rect 2550 330 2740 480
rect 2740 330 2820 480
rect 2550 320 2820 330
rect 30 -240 3240 -200
rect 30 -310 90 -240
rect 90 -310 3190 -240
rect 3190 -310 3240 -240
rect 30 -450 3240 -310
<< metal3 >>
rect -1218 1120 3368 1164
rect -1218 850 20 1120
rect 3250 850 3368 1120
rect -1218 840 3368 850
rect 60 690 730 760
rect 60 470 450 690
rect 720 470 730 690
rect 60 450 730 470
rect 790 690 2990 700
rect 790 620 810 690
rect 920 620 1840 690
rect 1950 620 2870 690
rect 2980 620 2990 690
rect 790 610 2990 620
rect 790 450 2450 610
rect 2540 490 3210 550
rect 280 380 2480 390
rect 280 310 290 380
rect 400 310 1320 380
rect 1430 310 2360 380
rect 2470 310 2480 380
rect 280 300 2480 310
rect 820 140 2480 300
rect 2540 320 2550 490
rect 2820 320 3210 490
rect 2540 160 3210 320
rect -1218 -200 3368 -170
rect -1218 -450 30 -200
rect 3240 -450 3368 -200
rect -1218 -568 3368 -450
<< labels >>
flabel metal3 2820 160 3210 550 0 FreeSans 800 0 0 0 INn
port 5 nsew
flabel metal3 790 450 2450 700 0 FreeSans 800 0 0 0 OUT
port 1 nsew
flabel metal3 30 -450 3240 -200 0 FreeSans 800 0 0 0 VSS
port 2 nsew
flabel metal3 20 850 3250 1120 0 FreeSans 800 0 0 0 VDD
port 3 nsew
flabel metal3 60 450 450 760 0 FreeSans 800 0 0 0 INp
port 4 nsew
flabel metal2 -480 -170 -40 110 0 FreeSans 1600 0 0 0 R
port 6 nsew
<< end >>
