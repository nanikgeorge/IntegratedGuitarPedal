magic
tech sky130A
magscale 1 2
timestamp 1713320270
<< nwell >>
rect -194 -164 194 198
<< pmos >>
rect -100 -64 100 136
<< pdiff >>
rect -158 124 -100 136
rect -158 -52 -146 124
rect -112 -52 -100 124
rect -158 -64 -100 -52
rect 100 124 158 136
rect 100 -52 112 124
rect 146 -52 158 124
rect 100 -64 158 -52
<< pdiffc >>
rect -146 -52 -112 124
rect 112 -52 146 124
<< poly >>
rect -100 136 100 162
rect -100 -111 100 -64
rect -100 -145 -84 -111
rect 84 -145 100 -111
rect -100 -161 100 -145
<< polycont >>
rect -84 -145 84 -111
<< locali >>
rect -146 124 -112 140
rect -146 -68 -112 -52
rect 112 124 146 140
rect 112 -68 146 -52
rect -100 -145 -84 -111
rect 84 -145 100 -111
<< viali >>
rect -146 -52 -112 124
rect 112 -52 146 124
rect -84 -145 84 -111
<< metal1 >>
rect -152 124 -106 136
rect -152 -52 -146 124
rect -112 -52 -106 124
rect -152 -64 -106 -52
rect 106 124 152 136
rect 106 -52 112 124
rect 146 -52 152 124
rect 106 -64 152 -52
rect -96 -111 96 -105
rect -96 -145 -84 -111
rect 84 -145 96 -111
rect -96 -151 96 -145
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 1 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
