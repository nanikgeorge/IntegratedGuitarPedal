* NGSPICE file created from opamp_flat.ext - technology: sky130A

.subckt myOpamp VDD OUT INp INn VSS
X0 a_320_185# VSS.t21 VSS.t22 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1 OUT.t6 INn.t0 a_578_185# VSS.t24 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2 VSS.t20 VSS.t18 VSS.t20 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X3 a_320_185# INp.t0 a_578_185# VSS.t26 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X4 VSS.t17 VSS.t14 VSS.t16 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0 ps=0 w=0.42 l=1
X5 VDD a_n476_n270# VSS sky130_fd_pr__res_xhigh_po_0p35 l=26.11
X6 a_320_185# a_320_185# VDD.t25 VDD.t24 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X7 a_578_185# a_n476_n270# VSS.t35 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X8 VSS.t13 VSS.t12 OUT.t1 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X9 VSS.t33 a_n476_n270# a_n476_n270# VSS.t24 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X10 VSS.t32 a_n476_n270# a_578_185# VSS.t23 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X11 a_n476_n270# a_n476_n270# VSS.t31 VSS.t30 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X12 VDD.t23 a_320_185# OUT.t10 VDD.t22 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X13 VDD.t21 a_320_185# a_320_185# VDD.t20 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X14 a_578_185# a_n476_n270# VSS.t29 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X15 VDD.t19 a_320_185# OUT.t8 VDD.t18 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X16 OUT.t5 INn.t1 a_578_185# VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X17 a_320_185# VDD.t3 VDD.t5 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X18 OUT.t7 a_320_185# VDD.t17 VDD.t16 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X19 a_320_185# a_320_185# VDD.t15 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X20 a_578_185# INp.t1 a_320_185# VSS.t30 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X21 VDD.t2 VDD.t0 OUT.t0 VDD.t1 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X22 a_578_185# INp.t2 a_320_185# VSS.t19 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X23 OUT.t4 INn.t2 a_578_185# VSS.t7 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X24 VSS.t11 VSS.t9 VSS.t11 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X25 VSS.t8 VSS.t6 VSS.t8 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X26 VSS.t27 a_n476_n270# a_578_185# VSS.t26 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X27 VSS.t5 VSS.t3 VSS.t5 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X28 a_320_185# INp.t3 a_578_185# VSS.t23 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X29 VDD.t26 a_n476_n270# VSS.t25 sky130_fd_pr__res_xhigh_po_0p35 l=0.16
X30 OUT.t11 a_320_185# VDD.t13 VDD.t12 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X31 a_578_185# INn.t3 OUT.t3 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X32 a_578_185# INp.t4 a_320_185# VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X33 VDD.t11 a_320_185# a_320_185# VDD.t10 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X34 a_578_185# INn.t4 OUT.t2 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X35 VDD.t9 a_320_185# a_320_185# VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X36 OUT.t9 a_320_185# VDD.t7 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X37 VSS.t2 VSS.t0 VSS.t2 VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
R0 VSS.n43 VSS.n36 27500
R1 VSS.t25 VSS.n43 10325.8
R2 VSS.n45 VSS.n18 10285.8
R3 VSS.n42 VSS.n18 10253
R4 VSS.n45 VSS.n19 10250
R5 VSS.n42 VSS.n19 10187.3
R6 VSS.n36 VSS.t10 1302.55
R7 VSS.t10 VSS.t7 803.966
R8 VSS.t7 VSS.t4 803.966
R9 VSS.t4 VSS.t26 803.966
R10 VSS.t26 VSS.t34 803.966
R11 VSS.t34 VSS.t24 803.966
R12 VSS.t30 VSS.t23 803.966
R13 VSS.t28 VSS.t1 803.966
R14 VSS.t1 VSS.t19 803.966
R15 VSS.t19 VSS.t15 803.966
R16 VSS.n47 VSS.n16 666.376
R17 VSS.n46 VSS.n17 665.019
R18 VSS.n39 VSS.n37 664.242
R19 VSS.n41 VSS.n40 661.915
R20 VSS.t15 VSS.t25 660.674
R21 VSS.n44 VSS.t23 629.462
R22 VSS.t24 VSS.n35 414.449
R23 VSS.n35 VSS.t30 389.519
R24 VSS.n26 VSS.t17 236.113
R25 VSS.t11 VSS.n3 235.764
R26 VSS.n31 VSS.n30 194.805
R27 VSS.n10 VSS.n9 194.542
R28 VSS.n33 VSS.n32 194.463
R29 VSS.n12 VSS.n11 194.463
R30 VSS.n27 VSS.n26 194.3
R31 VSS.n29 VSS.n28 194.3
R32 VSS.n8 VSS.n7 194.3
R33 VSS.n5 VSS.n4 194.3
R34 VSS.n36 VSS.n18 189.166
R35 VSS.n44 VSS.t28 174.505
R36 VSS.n23 VSS.t21 118.005
R37 VSS.n2 VSS.t12 118.005
R38 VSS.n24 VSS.t14 104.028
R39 VSS.n22 VSS.t18 104.028
R40 VSS.n21 VSS.t0 104.028
R41 VSS.n0 VSS.t3 104.028
R42 VSS.n6 VSS.t6 104.028
R43 VSS.n1 VSS.t9 104.028
R44 VSS.n23 VSS.t22 87.6949
R45 VSS.n2 VSS.t13 87.5315
R46 VSS.t25 VSS.n19 77.0353
R47 VSS.n30 VSS.t29 41.4291
R48 VSS.n30 VSS.t2 41.4291
R49 VSS.t20 VSS.n27 41.4291
R50 VSS.n27 VSS.t16 41.4291
R51 VSS.t2 VSS.n29 41.4291
R52 VSS.n29 VSS.t20 41.4291
R53 VSS.n32 VSS.t31 41.4291
R54 VSS.n32 VSS.t32 41.4291
R55 VSS.n9 VSS.t5 41.4291
R56 VSS.n9 VSS.t27 41.4291
R57 VSS.n8 VSS.t8 41.4291
R58 VSS.t5 VSS.n8 41.4291
R59 VSS.n4 VSS.t11 41.4291
R60 VSS.n4 VSS.t8 41.4291
R61 VSS.n11 VSS.t35 41.4291
R62 VSS.n11 VSS.t33 41.4291
R63 VSS.n35 VSS.n34 26.2219
R64 VSS.n40 VSS.n19 20.8934
R65 VSS.n37 VSS.n18 20.8934
R66 VSS.n42 VSS.n41 8.23994
R67 VSS.n43 VSS.n42 8.23994
R68 VSS.n46 VSS.n45 8.23994
R69 VSS.n45 VSS.n44 8.23994
R70 VSS.n38 VSS.n15 2.09737
R71 VSS.n48 VSS.n15 2.09737
R72 VSS.n38 VSS.n14 2.09113
R73 VSS.n41 VSS.n39 1.93989
R74 VSS.n49 VSS.n14 1.72862
R75 VSS.n40 VSS.n17 0.970197
R76 VSS.n47 VSS.n46 0.970197
R77 VSS.n37 VSS.n16 0.970197
R78 VSS.n33 VSS.n31 0.927299
R79 VSS.n12 VSS.n10 0.690273
R80 VSS.n31 VSS.n20 0.60675
R81 VSS.n31 VSS.n25 0.516045
R82 VSS.n21 VSS.n20 0.454213
R83 VSS.n49 VSS.n48 0.363
R84 VSS.n28 VSS.n20 0.347226
R85 VSS.n16 VSS.n14 0.344944
R86 VSS.n17 VSS.n15 0.344944
R87 VSS.n22 VSS.n21 0.319807
R88 VSS.n25 VSS.n24 0.291342
R89 VSS.n28 VSS.n25 0.22669
R90 VSS.n13 VSS.n12 0.216409
R91 VSS.n34 VSS.n33 0.210727
R92 VSS.n26 VSS.n25 0.158238
R93 VSS.n39 VSS.n38 0.135283
R94 VSS.n48 VSS.n47 0.135283
R95 VSS VSS.n50 0.11003
R96 VSS.n50 VSS.n13 0.0961731
R97 VSS.n24 VSS.n23 0.0714406
R98 VSS.n50 VSS.n49 0.0599231
R99 VSS.n5 VSS.n1 0.0429342
R100 VSS.n6 VSS.n5 0.0429342
R101 VSS.n7 VSS.n6 0.0429342
R102 VSS.n7 VSS.n0 0.0429342
R103 VSS.n3 VSS.n2 0.0389615
R104 VSS.n10 VSS.n0 0.0340526
R105 VSS.n25 VSS.n22 0.0289653
R106 VSS.n3 VSS.n1 0.00773684
R107 VSS.n34 VSS.n13 0.00618182
R108 INn.n0 INn.t1 118.769
R109 INn.n3 INn.t2 118.005
R110 INn.n2 INn.t3 118.005
R111 INn.n1 INn.t0 118.005
R112 INn.n0 INn.t4 118.005
R113 INn INn.n3 3.33334
R114 INn.n1 INn.n0 2.66195
R115 INn.n3 INn.n2 2.55325
R116 INn.n2 INn.n1 0.764886
R117 OUT.n9 OUT.n7 204.206
R118 OUT.n5 OUT.n3 204.206
R119 OUT.n2 OUT.n0 204.206
R120 OUT.n9 OUT.n8 71.1729
R121 OUT.n5 OUT.n4 71.1729
R122 OUT.n2 OUT.n1 71.1729
R123 OUT.n7 OUT.t8 28.5655
R124 OUT.n7 OUT.t11 28.5655
R125 OUT.n3 OUT.t10 28.5655
R126 OUT.n3 OUT.t7 28.5655
R127 OUT.n0 OUT.t0 28.5655
R128 OUT.n0 OUT.t9 28.5655
R129 OUT.n8 OUT.t2 17.4005
R130 OUT.n8 OUT.t5 17.4005
R131 OUT.n4 OUT.t3 17.4005
R132 OUT.n4 OUT.t6 17.4005
R133 OUT.n1 OUT.t1 17.4005
R134 OUT.n1 OUT.t4 17.4005
R135 OUT.n6 OUT.n2 3.7629
R136 OUT.n6 OUT.n5 3.4105
R137 OUT.n10 OUT.n9 3.4105
R138 OUT.n10 OUT.n6 0.19414
R139 OUT OUT.n10 0.0146
R140 INp.n0 INp.t4 118.769
R141 INp.n3 INp.t2 118.621
R142 INp.n2 INp.t3 118.005
R143 INp.n1 INp.t1 118.005
R144 INp.n0 INp.t0 118.005
R145 INp INp.n3 2.77717
R146 INp.n1 INp.n0 2.66195
R147 INp.n3 INp.n2 1.71868
R148 INp.n2 INp.n1 0.764886
R149 VDD.n14 VDD.n13 18810
R150 VDD.n15 VDD.n14 18786.2
R151 VDD.n15 VDD.n6 18786.2
R152 VDD.n13 VDD.n6 18667.5
R153 VDD.n16 VDD.n4 7334.54
R154 VDD.n12 VDD.n5 7332.73
R155 VDD.n16 VDD.n5 7312.73
R156 VDD.n12 VDD.n4 7300
R157 VDD.n10 VDD.n8 781.188
R158 VDD.n18 VDD.n2 779.442
R159 VDD.n17 VDD.n3 779.056
R160 VDD.n11 VDD.n7 778.668
R161 VDD.t6 VDD.t1 478.712
R162 VDD.t20 VDD.t6 478.712
R163 VDD.t14 VDD.t20 478.712
R164 VDD.t22 VDD.t14 478.712
R165 VDD.t16 VDD.t22 478.712
R166 VDD.t10 VDD.t24 478.712
R167 VDD.t24 VDD.t18 478.712
R168 VDD.t18 VDD.t12 478.712
R169 VDD.t12 VDD.t8 478.712
R170 VDD.t8 VDD.t4 478.712
R171 VDD.n31 VDD.t10 269.043
R172 VDD.n32 VDD.t26 264.031
R173 VDD.n26 VDD.t5 228.215
R174 VDD.n21 VDD.t2 228.215
R175 VDD.n31 VDD.t16 209.668
R176 VDD.n28 VDD.n27 199.851
R177 VDD.n30 VDD.n29 199.851
R178 VDD.n23 VDD.n22 199.851
R179 VDD.n25 VDD.n24 199.851
R180 VDD.n35 VDD.n34 199.851
R181 VDD.n21 VDD.t0 120.855
R182 VDD.n26 VDD.t3 120.749
R183 VDD.n32 VDD.n31 38.8096
R184 VDD.n27 VDD.t13 28.5655
R185 VDD.n27 VDD.t9 28.5655
R186 VDD.n29 VDD.t25 28.5655
R187 VDD.n29 VDD.t19 28.5655
R188 VDD.n22 VDD.t7 28.5655
R189 VDD.n22 VDD.t21 28.5655
R190 VDD.n24 VDD.t15 28.5655
R191 VDD.n24 VDD.t23 28.5655
R192 VDD.n34 VDD.t17 28.5655
R193 VDD.n34 VDD.t11 28.5655
R194 VDD.n8 VDD.n5 5.0005
R195 VDD.n14 VDD.n5 5.0005
R196 VDD.n7 VDD.n4 4.86892
R197 VDD.n6 VDD.n4 4.86892
R198 VDD.n19 VDD.n1 2.4755
R199 VDD.n9 VDD.n1 2.4755
R200 VDD.n9 VDD.n0 2.463
R201 VDD.n17 VDD.n16 2.34227
R202 VDD.n16 VDD.n15 2.34227
R203 VDD.n12 VDD.n11 2.34227
R204 VDD.n13 VDD.n12 2.34227
R205 VDD.n20 VDD.n0 2.10363
R206 VDD.n18 VDD.n17 1.93989
R207 VDD.n7 VDD.n2 0.970197
R208 VDD.n11 VDD.n10 0.970197
R209 VDD.n8 VDD.n3 0.970197
R210 VDD.n23 VDD.n21 0.890989
R211 VDD.n28 VDD.n26 0.760446
R212 VDD.n30 VDD.n28 0.40675
R213 VDD.n25 VDD.n23 0.40675
R214 VDD.n35 VDD.n25 0.40675
R215 VDD.n20 VDD.n19 0.359875
R216 VDD.n3 VDD.n1 0.258833
R217 VDD.n2 VDD.n0 0.258833
R218 VDD.n35 VDD.n33 0.208833
R219 VDD.n33 VDD.n30 0.188
R220 VDD.n33 VDD.n32 0.1865
R221 VDD.n10 VDD.n9 0.121279
R222 VDD.n19 VDD.n18 0.121279
R223 VDD VDD.n36 0.117178
R224 VDD.n36 VDD.n35 0.0948367
R225 VDD.n36 VDD.n20 0.0691538
C0 OUT INn 1.03193f
C1 VDD INn 0.172037f
C2 a_320_185# OUT 2.35058f
C3 OUT a_n476_n270# 0.001336f
C4 a_320_185# VDD 4.40463f
C5 VDD a_n476_n270# 0.09688f
C6 OUT INp 0.763432f
C7 VDD INp 0.673697f
C8 a_578_185# OUT 0.662032f
C9 VDD a_578_185# 0.137313f
C10 a_320_185# INn 0.849481f
C11 a_n476_n270# INn 1.1307f
C12 a_320_185# a_n476_n270# 0.27522f
C13 INp INn 0.500623f
C14 a_320_185# INp 3.09291f
C15 a_n476_n270# INp 0.162656f
C16 a_578_185# INn 1.23455f
C17 a_320_185# a_578_185# 1.57848f
C18 a_578_185# a_n476_n270# 1.5318f
C19 a_578_185# INp 0.763261f
C20 VDD OUT 1.99539f
C21 INn VSS 2.51255f
C22 INp VSS 3.09822f
C23 OUT VSS 0.502824f
C24 VDD VSS 41.529198f
C25 a_n476_n270# VSS 5.4076f
C26 a_578_185# VSS 1.59044f
C27 a_320_185# VSS 2.69418f
C28 VDD.n0 VSS 0.175287f
C29 VDD.n1 VSS 0.189777f
C30 VDD.n2 VSS 0.03108f
C31 VDD.n3 VSS 0.031065f
C32 VDD.n4 VSS 0.062168f
C33 VDD.n5 VSS 0.062214f
C34 VDD.n6 VSS 0.188955f
C35 VDD.n7 VSS 0.03105f
C36 VDD.n8 VSS 0.031149f
C37 VDD.n9 VSS 0.185674f
C38 VDD.n10 VSS 0.030967f
C39 VDD.n11 VSS 0.030868f
C40 VDD.n12 VSS 0.061797f
C41 VDD.n13 VSS 0.185434f
C42 VDD.n14 VSS 0.18966f
C43 VDD.n15 VSS 0.185914f
C44 VDD.n16 VSS 0.061858f
C45 VDD.n17 VSS 0.030921f
C46 VDD.n18 VSS 0.030937f
C47 VDD.n19 VSS 0.106374f
C48 VDD.n20 VSS 0.198469f
C49 VDD.t0 VSS 0.010891f
C50 VDD.t2 VSS 0.002466f
C51 VDD.n21 VSS 0.014271f
C52 VDD.t7 VSS 6.71e-19
C53 VDD.t21 VSS 6.71e-19
C54 VDD.n22 VSS 0.001388f
C55 VDD.n23 VSS 0.027564f
C56 VDD.t15 VSS 6.71e-19
C57 VDD.t23 VSS 6.71e-19
C58 VDD.n24 VSS 0.001388f
C59 VDD.n25 VSS 0.023172f
C60 VDD.t3 VSS 0.010883f
C61 VDD.t5 VSS 0.002466f
C62 VDD.n26 VSS 0.024709f
C63 VDD.t13 VSS 6.71e-19
C64 VDD.t9 VSS 6.71e-19
C65 VDD.n27 VSS 0.001388f
C66 VDD.n28 VSS 0.033097f
C67 VDD.t25 VSS 6.71e-19
C68 VDD.t19 VSS 6.71e-19
C69 VDD.n29 VSS 0.001388f
C70 VDD.n30 VSS 0.020255f
C71 VDD.t1 VSS 0.03828f
C72 VDD.t6 VSS 0.030576f
C73 VDD.t20 VSS 0.030576f
C74 VDD.t14 VSS 0.030576f
C75 VDD.t22 VSS 0.030576f
C76 VDD.t16 VSS 0.021984f
C77 VDD.t4 VSS 0.03828f
C78 VDD.t8 VSS 0.030576f
C79 VDD.t12 VSS 0.030576f
C80 VDD.t18 VSS 0.030576f
C81 VDD.t24 VSS 0.030576f
C82 VDD.t10 VSS 0.02388f
C83 VDD.n31 VSS -0.017931f
C84 VDD.t26 VSS 0.025145f
C85 VDD.n32 VSS 0.038891f
C86 VDD.n33 VSS 0.005278f
C87 VDD.t17 VSS 6.71e-19
C88 VDD.t11 VSS 6.71e-19
C89 VDD.n34 VSS 0.001388f
C90 VDD.n35 VSS 0.022776f
C91 VDD.n36 VSS 1.00176f
C92 INp.t4 VSS 0.192033f
C93 INp.t0 VSS 0.191404f
C94 INp.n0 VSS 0.237081f
C95 INp.t1 VSS 0.191404f
C96 INp.n1 VSS 0.139872f
C97 INp.t3 VSS 0.191404f
C98 INp.n2 VSS 0.121401f
C99 INp.t2 VSS 0.191893f
C100 INp.n3 VSS 0.332858f
C101 OUT.t0 VSS 0.007912f
C102 OUT.t9 VSS 0.007912f
C103 OUT.n0 VSS 0.018165f
C104 OUT.t1 VSS 0.007912f
C105 OUT.t4 VSS 0.007912f
C106 OUT.n1 VSS 0.023194f
C107 OUT.n2 VSS 0.320387f
C108 OUT.t10 VSS 0.007912f
C109 OUT.t7 VSS 0.007912f
C110 OUT.n3 VSS 0.018165f
C111 OUT.t3 VSS 0.007912f
C112 OUT.t6 VSS 0.007912f
C113 OUT.n4 VSS 0.023194f
C114 OUT.n5 VSS 0.306564f
C115 OUT.n6 VSS 0.848589f
C116 OUT.t8 VSS 0.007912f
C117 OUT.t11 VSS 0.007912f
C118 OUT.n7 VSS 0.018164f
C119 OUT.t2 VSS 0.007912f
C120 OUT.t5 VSS 0.007912f
C121 OUT.n8 VSS 0.023194f
C122 OUT.n9 VSS 0.303018f
C123 OUT.n10 VSS 0.376845f
.ends

