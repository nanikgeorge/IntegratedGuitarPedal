magic
tech sky130A
magscale 1 2
timestamp 1713319136
<< error_p >>
rect 524 100 610 132
rect 646 96 768 264
rect 560 64 768 96
rect 600 0 768 64
<< nwell >>
rect -20 1120 660 1380
rect 0 96 646 1120
rect 0 0 560 96
rect 600 0 646 96
<< nmos >>
rect 94 -1087 294 -87
rect 352 -1087 552 -87
<< pmos >>
rect 94 100 294 1100
rect 352 100 552 1100
<< ndiff >>
rect 36 -99 94 -87
rect 36 -1075 48 -99
rect 82 -1075 94 -99
rect 36 -1087 94 -1075
rect 294 -99 352 -87
rect 294 -1075 306 -99
rect 340 -1075 352 -99
rect 294 -1087 352 -1075
rect 552 -99 610 -87
rect 552 -1075 564 -99
rect 598 -1075 610 -99
rect 552 -1087 610 -1075
<< pdiff >>
rect 36 1088 94 1100
rect 36 112 48 1088
rect 82 112 94 1088
rect 36 100 94 112
rect 294 1088 352 1100
rect 294 112 306 1088
rect 340 112 352 1088
rect 294 100 352 112
rect 552 1088 610 1100
rect 552 112 564 1088
rect 598 112 610 1088
rect 552 100 610 112
<< ndiffc >>
rect 48 -1075 82 -99
rect 306 -1075 340 -99
rect 564 -1075 598 -99
<< pdiffc >>
rect 48 112 82 1088
rect 306 112 340 1088
rect 564 112 598 1088
<< psubdiff >>
rect 750 -130 1072 -106
rect 750 -1074 1072 -1050
<< nsubdiff >>
rect 40 1300 600 1340
rect 40 1200 80 1300
rect 560 1200 600 1300
rect 40 1160 600 1200
<< psubdiffcont >>
rect 750 -1050 1072 -130
<< nsubdiffcont >>
rect 80 1200 560 1300
<< poly >>
rect 94 1100 294 1126
rect 352 1100 552 1126
rect 94 53 294 100
rect 94 19 110 53
rect 278 19 294 53
rect 94 3 294 19
rect 352 53 552 100
rect 352 19 368 53
rect 536 19 552 53
rect 352 3 552 19
rect 94 -87 294 -61
rect 352 -87 552 -61
rect 94 -1125 294 -1087
rect 94 -1159 110 -1125
rect 278 -1159 294 -1125
rect 94 -1175 294 -1159
rect 352 -1125 552 -1087
rect 352 -1159 368 -1125
rect 536 -1159 552 -1125
rect 352 -1175 552 -1159
<< polycont >>
rect 110 19 278 53
rect 368 19 536 53
rect 110 -1159 278 -1125
rect 368 -1159 536 -1125
<< locali >>
rect 60 1300 580 1320
rect 60 1200 80 1300
rect 560 1200 580 1300
rect 60 1180 580 1200
rect 48 1088 82 1104
rect 48 96 82 112
rect 306 1088 340 1104
rect 306 96 340 112
rect 564 1088 598 1104
rect 564 96 598 112
rect 94 19 110 53
rect 278 19 294 53
rect 352 19 368 53
rect 536 19 552 53
rect 48 -99 82 -83
rect 48 -1091 82 -1075
rect 306 -99 340 -83
rect 306 -1091 340 -1075
rect 564 -99 598 -83
rect 750 -130 1072 -114
rect 750 -1066 1072 -1050
rect 564 -1091 598 -1075
rect 94 -1159 110 -1125
rect 278 -1159 294 -1125
rect 352 -1159 368 -1125
rect 536 -1159 552 -1125
<< viali >>
rect 80 1200 560 1300
rect 48 112 82 1088
rect 306 112 340 1088
rect 564 112 598 1088
rect 110 19 278 53
rect 368 19 536 53
rect 48 -1075 82 -99
rect 306 -1075 340 -99
rect 564 -1075 598 -99
rect 820 -1040 980 -140
rect 110 -1159 278 -1125
rect 368 -1159 536 -1125
<< metal1 >>
rect 40 1300 600 1340
rect 40 1200 80 1300
rect 560 1200 600 1300
rect 40 1160 600 1200
rect 38 1100 80 1120
rect 38 1088 88 1100
rect 38 112 48 1088
rect 82 112 88 1088
rect 38 100 88 112
rect 280 1088 360 1160
rect 280 112 306 1088
rect 340 112 360 1088
rect 280 100 360 112
rect 558 1088 682 1100
rect 558 112 564 1088
rect 598 112 682 1088
rect 558 100 682 112
rect 38 60 80 100
rect 580 96 682 100
rect 38 53 560 60
rect 38 19 110 53
rect 278 19 368 53
rect 536 19 560 53
rect 38 -20 560 19
rect 38 -22 302 -20
rect 38 -87 80 -22
rect 600 -80 682 96
rect 580 -87 682 -80
rect 38 -99 88 -87
rect 38 -1075 48 -99
rect 82 -1075 88 -99
rect 300 -99 346 -87
rect 300 -220 306 -99
rect 220 -980 306 -220
rect 38 -1080 88 -1075
rect 42 -1087 88 -1080
rect 300 -1075 306 -980
rect 340 -220 346 -99
rect 558 -99 682 -87
rect 340 -980 420 -220
rect 340 -1075 346 -980
rect 300 -1087 346 -1075
rect 558 -1075 564 -99
rect 598 -1075 682 -99
rect 558 -1080 682 -1075
rect 744 -140 1116 -18
rect 744 -1040 820 -140
rect 980 -1040 1116 -140
rect 558 -1087 604 -1080
rect 98 -1120 290 -1119
rect 356 -1120 548 -1119
rect 80 -1125 300 -1120
rect 80 -1159 110 -1125
rect 278 -1159 300 -1125
rect 80 -1280 300 -1159
rect 340 -1125 560 -1120
rect 340 -1159 368 -1125
rect 536 -1159 560 -1125
rect 340 -1280 560 -1159
rect 744 -1168 1116 -1040
<< labels >>
flabel metal1 220 -980 420 -220 0 FreeSans 160 0 0 0 currentOut
port 5 nsew
flabel metal1 744 -1168 1116 -18 0 FreeSans 160 0 0 0 VSS
port 6 nsew
flabel metal1 280 100 360 1200 0 FreeSans 160 0 0 0 VDD
port 2 nsew
flabel metal1 80 -1280 300 -1120 0 FreeSans 160 0 0 0 inp
port 3 nsew
flabel metal1 340 -1280 560 -1120 0 FreeSans 160 0 0 0 inn
port 4 nsew
<< end >>
