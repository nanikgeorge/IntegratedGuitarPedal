* NGSPICE file created from tt_um_flat.ext - technology: sky130A

.subckt myOpamp OUT VSS VDD INp INn
X0 a_320_185# VSS.t22 VSS.t23 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1 OUT.t4 INn.t0 a_578_185# VSS.t33 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2 VSS.t21 VSS.t20 VSS.t21 VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0 ps=0 w=0.5 l=1
X3 a_320_185# INp.t0 a_578_185# VSS.t26 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X4 VSS.t19 VSS.t16 VSS.t18 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=1
X5 VDD a_n476_n270# VSS sky130_fd_pr__res_xhigh_po_0p35 l=26.11
X6 a_320_185# a_320_185# VDD.t19 VDD.t18 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X7 a_578_185# a_n476_n270# VSS.t35 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=1
X8 VSS.t15 VSS.t14 OUT.t10 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X9 VSS.t34 a_n476_n270# a_n476_n270# VSS.t33 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=1
X10 VSS.t32 a_n476_n270# a_578_185# VSS.t31 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=1
X11 a_n476_n270# a_n476_n270# VSS.t30 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=1
X12 VDD.t17 a_320_185# OUT.t7 VDD.t16 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X13 VDD.t15 a_320_185# a_320_185# VDD.t14 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X14 a_578_185# a_n476_n270# VSS.t28 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=1
X15 VDD.t13 a_320_185# OUT.t8 VDD.t12 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X16 OUT.t3 INn.t1 a_578_185# VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X17 a_320_185# VDD.t24 VDD.t26 VDD.t25 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X18 OUT.t5 a_320_185# VDD.t11 VDD.t10 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X19 a_320_185# a_320_185# VDD.t9 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X20 a_578_185# INp.t1 a_320_185# VSS.t29 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X21 VDD.t23 VDD.t21 OUT.t11 VDD.t22 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X22 a_578_185# INp.t2 a_320_185# VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X23 OUT.t2 INn.t2 a_578_185# VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X24 VSS.t13 VSS.t11 VSS.t13 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0 ps=0 w=0.5 l=1
X25 VSS.t10 VSS.t9 VSS.t10 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0 ps=0 w=0.5 l=1
X26 VSS.t27 a_n476_n270# a_578_185# VSS.t26 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=1
X27 VSS.t8 VSS.t6 VSS.t8 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0 ps=0 w=0.5 l=1
X28 a_320_185# INp.t3 a_578_185# VSS.t31 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X29 VDD.t20 a_n476_n270# VSS.t24 sky130_fd_pr__res_xhigh_po_0p35 l=0.16
X30 OUT.t6 a_320_185# VDD.t7 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X31 a_578_185# INn.t3 OUT.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X32 a_578_185# INp.t4 a_320_185# VSS.t7 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X33 VDD.t5 a_320_185# a_320_185# VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X34 a_578_185# INn.t4 OUT.t0 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X35 VDD.t3 a_320_185# a_320_185# VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X36 OUT.t9 a_320_185# VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X37 VSS.t5 VSS.t3 VSS.t5 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0 ps=0 w=0.5 l=1
R0 VSS.n42 VSS.n35 27500
R1 VSS.t24 VSS.n42 10325.8
R2 VSS.n44 VSS.n18 10285.8
R3 VSS.n41 VSS.n18 10253
R4 VSS.n44 VSS.n19 10250
R5 VSS.n41 VSS.n19 10187.3
R6 VSS.n35 VSS.t12 1302.55
R7 VSS.t12 VSS.t2 803.966
R8 VSS.t2 VSS.t7 803.966
R9 VSS.t7 VSS.t26 803.966
R10 VSS.t26 VSS.t0 803.966
R11 VSS.t0 VSS.t33 803.966
R12 VSS.t29 VSS.t31 803.966
R13 VSS.t25 VSS.t4 803.966
R14 VSS.t4 VSS.t1 803.966
R15 VSS.t1 VSS.t17 803.966
R16 VSS.n46 VSS.n16 666.376
R17 VSS.n45 VSS.n17 665.019
R18 VSS.n38 VSS.n36 664.242
R19 VSS.n40 VSS.n39 661.915
R20 VSS.t17 VSS.t24 660.674
R21 VSS.n43 VSS.t31 629.462
R22 VSS.t33 VSS.n34 414.449
R23 VSS.n34 VSS.t29 389.519
R24 VSS.t13 VSS.n3 229.136
R25 VSS.n22 VSS.t19 229.135
R26 VSS.n30 VSS.n29 194.571
R27 VSS.n10 VSS.n9 194.538
R28 VSS.n32 VSS.n31 194.47
R29 VSS.n12 VSS.n11 194.47
R30 VSS.n25 VSS.n24 194.3
R31 VSS.n28 VSS.n27 194.3
R32 VSS.n8 VSS.n7 194.3
R33 VSS.n5 VSS.n4 194.3
R34 VSS.n35 VSS.n18 189.166
R35 VSS.n43 VSS.t25 174.505
R36 VSS.n21 VSS.t22 118.005
R37 VSS.n2 VSS.t14 118.005
R38 VSS.n23 VSS.t16 105.956
R39 VSS.n26 VSS.t20 105.956
R40 VSS.n20 VSS.t3 105.956
R41 VSS.n0 VSS.t6 105.956
R42 VSS.n6 VSS.t9 105.956
R43 VSS.n1 VSS.t11 105.956
R44 VSS.n21 VSS.t23 87.6949
R45 VSS.n2 VSS.t15 87.5315
R46 VSS.t24 VSS.n19 77.0353
R47 VSS.n29 VSS.t28 34.8005
R48 VSS.n29 VSS.t5 34.8005
R49 VSS.n24 VSS.t21 34.8005
R50 VSS.n24 VSS.t18 34.8005
R51 VSS.t5 VSS.n28 34.8005
R52 VSS.n28 VSS.t21 34.8005
R53 VSS.n31 VSS.t30 34.8005
R54 VSS.n31 VSS.t32 34.8005
R55 VSS.n9 VSS.t8 34.8005
R56 VSS.n9 VSS.t27 34.8005
R57 VSS.n8 VSS.t10 34.8005
R58 VSS.t8 VSS.n8 34.8005
R59 VSS.n4 VSS.t13 34.8005
R60 VSS.n4 VSS.t10 34.8005
R61 VSS.n11 VSS.t35 34.8005
R62 VSS.n11 VSS.t34 34.8005
R63 VSS.n34 VSS.n33 26.2219
R64 VSS.n39 VSS.n19 20.8934
R65 VSS.n36 VSS.n18 20.8934
R66 VSS.n41 VSS.n40 8.23994
R67 VSS.n42 VSS.n41 8.23994
R68 VSS.n45 VSS.n44 8.23994
R69 VSS.n44 VSS.n43 8.23994
R70 VSS.n37 VSS.n15 2.09737
R71 VSS.n47 VSS.n15 2.09737
R72 VSS.n37 VSS.n14 2.09113
R73 VSS.n40 VSS.n38 1.93989
R74 VSS.n48 VSS.n14 1.72862
R75 VSS.n39 VSS.n17 0.970197
R76 VSS.n46 VSS.n45 0.970197
R77 VSS.n36 VSS.n16 0.970197
R78 VSS.n32 VSS.n30 0.754477
R79 VSS.n12 VSS.n10 0.715273
R80 VSS.n48 VSS.n47 0.363
R81 VSS.n16 VSS.n14 0.344944
R82 VSS.n17 VSS.n15 0.344944
R83 VSS.n13 VSS.n12 0.216409
R84 VSS.n33 VSS.n32 0.210727
R85 VSS.n38 VSS.n37 0.135283
R86 VSS.n47 VSS.n46 0.135283
R87 VSS VSS.n49 0.11003
R88 VSS.n49 VSS.n13 0.0961731
R89 VSS.n49 VSS.n48 0.0599231
R90 VSS.n27 VSS.n20 0.0429342
R91 VSS.n27 VSS.n26 0.0429342
R92 VSS.n26 VSS.n25 0.0429342
R93 VSS.n25 VSS.n23 0.0429342
R94 VSS.n5 VSS.n1 0.0429342
R95 VSS.n6 VSS.n5 0.0429342
R96 VSS.n7 VSS.n6 0.0429342
R97 VSS.n7 VSS.n0 0.0429342
R98 VSS.n22 VSS.n21 0.0405
R99 VSS.n3 VSS.n2 0.0389615
R100 VSS.n30 VSS.n20 0.0347105
R101 VSS.n10 VSS.n0 0.0340526
R102 VSS.n23 VSS.n22 0.00872368
R103 VSS.n3 VSS.n1 0.00773684
R104 VSS.n33 VSS.n13 0.00618182
R105 INn.n0 INn.t1 118.769
R106 INn.n3 INn.t2 118.005
R107 INn.n2 INn.t3 118.005
R108 INn.n1 INn.t0 118.005
R109 INn.n0 INn.t4 118.005
R110 INn INn.n3 3.33334
R111 INn.n1 INn.n0 2.66195
R112 INn.n3 INn.n2 2.55325
R113 INn.n2 INn.n1 0.764886
R114 OUT.n9 OUT.n7 204.206
R115 OUT.n5 OUT.n3 204.206
R116 OUT.n2 OUT.n0 204.206
R117 OUT.n9 OUT.n8 71.1729
R118 OUT.n5 OUT.n4 71.1729
R119 OUT.n2 OUT.n1 71.1729
R120 OUT.n7 OUT.t8 28.5655
R121 OUT.n7 OUT.t6 28.5655
R122 OUT.n3 OUT.t7 28.5655
R123 OUT.n3 OUT.t5 28.5655
R124 OUT.n0 OUT.t11 28.5655
R125 OUT.n0 OUT.t9 28.5655
R126 OUT.n8 OUT.t0 17.4005
R127 OUT.n8 OUT.t3 17.4005
R128 OUT.n4 OUT.t1 17.4005
R129 OUT.n4 OUT.t4 17.4005
R130 OUT.n1 OUT.t10 17.4005
R131 OUT.n1 OUT.t2 17.4005
R132 OUT.n6 OUT.n2 3.7629
R133 OUT.n6 OUT.n5 3.4105
R134 OUT.n10 OUT.n9 3.4105
R135 OUT.n10 OUT.n6 0.19414
R136 OUT OUT.n10 0.0146
R137 INp.n0 INp.t4 118.769
R138 INp.n3 INp.t2 118.621
R139 INp.n2 INp.t3 118.005
R140 INp.n1 INp.t1 118.005
R141 INp.n0 INp.t0 118.005
R142 INp INp.n3 2.77717
R143 INp.n1 INp.n0 2.66195
R144 INp.n3 INp.n2 1.71868
R145 INp.n2 INp.n1 0.764886
R146 VDD.n14 VDD.n13 18810
R147 VDD.n15 VDD.n14 18786.2
R148 VDD.n15 VDD.n6 18786.2
R149 VDD.n13 VDD.n6 18667.5
R150 VDD.n16 VDD.n4 7334.54
R151 VDD.n12 VDD.n5 7332.73
R152 VDD.n16 VDD.n5 7312.73
R153 VDD.n12 VDD.n4 7300
R154 VDD.n10 VDD.n8 781.188
R155 VDD.n18 VDD.n2 779.442
R156 VDD.n17 VDD.n3 779.056
R157 VDD.n11 VDD.n7 778.668
R158 VDD.t0 VDD.t22 478.712
R159 VDD.t14 VDD.t0 478.712
R160 VDD.t8 VDD.t14 478.712
R161 VDD.t16 VDD.t8 478.712
R162 VDD.t10 VDD.t16 478.712
R163 VDD.t4 VDD.t18 478.712
R164 VDD.t18 VDD.t12 478.712
R165 VDD.t12 VDD.t6 478.712
R166 VDD.t6 VDD.t2 478.712
R167 VDD.t2 VDD.t25 478.712
R168 VDD.n31 VDD.t4 269.043
R169 VDD.n32 VDD.t20 264.031
R170 VDD.n26 VDD.t26 228.215
R171 VDD.n21 VDD.t23 228.215
R172 VDD.n31 VDD.t10 209.668
R173 VDD.n28 VDD.n27 199.851
R174 VDD.n30 VDD.n29 199.851
R175 VDD.n23 VDD.n22 199.851
R176 VDD.n25 VDD.n24 199.851
R177 VDD.n35 VDD.n34 199.851
R178 VDD.n21 VDD.t21 120.855
R179 VDD.n26 VDD.t24 120.749
R180 VDD.n32 VDD.n31 38.8096
R181 VDD.n27 VDD.t7 28.5655
R182 VDD.n27 VDD.t3 28.5655
R183 VDD.n29 VDD.t19 28.5655
R184 VDD.n29 VDD.t13 28.5655
R185 VDD.n22 VDD.t1 28.5655
R186 VDD.n22 VDD.t15 28.5655
R187 VDD.n24 VDD.t9 28.5655
R188 VDD.n24 VDD.t17 28.5655
R189 VDD.n34 VDD.t11 28.5655
R190 VDD.n34 VDD.t5 28.5655
R191 VDD.n8 VDD.n5 5.0005
R192 VDD.n14 VDD.n5 5.0005
R193 VDD.n7 VDD.n4 4.86892
R194 VDD.n6 VDD.n4 4.86892
R195 VDD.n19 VDD.n1 2.4755
R196 VDD.n9 VDD.n1 2.4755
R197 VDD.n9 VDD.n0 2.463
R198 VDD.n17 VDD.n16 2.34227
R199 VDD.n16 VDD.n15 2.34227
R200 VDD.n12 VDD.n11 2.34227
R201 VDD.n13 VDD.n12 2.34227
R202 VDD.n20 VDD.n0 2.10363
R203 VDD.n18 VDD.n17 1.93989
R204 VDD.n7 VDD.n2 0.970197
R205 VDD.n11 VDD.n10 0.970197
R206 VDD.n8 VDD.n3 0.970197
R207 VDD.n23 VDD.n21 0.890989
R208 VDD.n28 VDD.n26 0.760446
R209 VDD.n30 VDD.n28 0.40675
R210 VDD.n25 VDD.n23 0.40675
R211 VDD.n35 VDD.n25 0.40675
R212 VDD.n20 VDD.n19 0.359875
R213 VDD.n3 VDD.n1 0.258833
R214 VDD.n2 VDD.n0 0.258833
R215 VDD.n35 VDD.n33 0.208833
R216 VDD.n33 VDD.n30 0.188
R217 VDD.n33 VDD.n32 0.1865
R218 VDD.n10 VDD.n9 0.121279
R219 VDD.n19 VDD.n18 0.121279
R220 VDD VDD.n36 0.117178
R221 VDD.n36 VDD.n35 0.0948367
R222 VDD.n36 VDD.n20 0.0691538
C0 INn OUT 1.03193f
C1 OUT a_n476_n270# 0.001186f
C2 INp OUT 0.763432f
C3 INn a_n476_n270# 1.22161f
C4 INp INn 0.500623f
C5 INp a_n476_n270# 0.1757f
C6 VDD a_578_185# 0.137337f
C7 VDD a_320_185# 4.40463f
C8 a_320_185# a_578_185# 1.57846f
C9 VDD OUT 1.99539f
C10 OUT a_578_185# 0.662059f
C11 a_320_185# OUT 2.35058f
C12 INn VDD 0.172037f
C13 VDD a_n476_n270# 0.096865f
C14 INn a_578_185# 1.23359f
C15 a_578_185# a_n476_n270# 1.482f
C16 INn a_320_185# 0.849481f
C17 INp VDD 0.673697f
C18 a_320_185# a_n476_n270# 0.272362f
C19 INp a_578_185# 0.763231f
C20 INp a_320_185# 3.09291f
C21 INn VSS 2.53371f
C22 INp VSS 3.09212f
C23 OUT VSS 0.503017f
C24 VDD VSS 41.529198f
C25 a_n476_n270# VSS 5.36992f
C26 a_578_185# VSS 1.63087f
C27 a_320_185# VSS 2.69798f
C28 VDD.n0 VSS 0.175287f
C29 VDD.n1 VSS 0.189777f
C30 VDD.n2 VSS 0.03108f
C31 VDD.n3 VSS 0.031065f
C32 VDD.n4 VSS 0.062168f
C33 VDD.n5 VSS 0.062214f
C34 VDD.n6 VSS 0.188955f
C35 VDD.n7 VSS 0.03105f
C36 VDD.n8 VSS 0.031149f
C37 VDD.n9 VSS 0.185674f
C38 VDD.n10 VSS 0.030967f
C39 VDD.n11 VSS 0.030868f
C40 VDD.n12 VSS 0.061797f
C41 VDD.n13 VSS 0.185434f
C42 VDD.n14 VSS 0.18966f
C43 VDD.n15 VSS 0.185914f
C44 VDD.n16 VSS 0.061858f
C45 VDD.n17 VSS 0.030921f
C46 VDD.n18 VSS 0.030937f
C47 VDD.n19 VSS 0.106374f
C48 VDD.n20 VSS 0.198469f
C49 VDD.t21 VSS 0.010891f
C50 VDD.t23 VSS 0.002466f
C51 VDD.n21 VSS 0.014271f
C52 VDD.t1 VSS 6.71e-19
C53 VDD.t15 VSS 6.71e-19
C54 VDD.n22 VSS 0.001388f
C55 VDD.n23 VSS 0.027564f
C56 VDD.t9 VSS 6.71e-19
C57 VDD.t17 VSS 6.71e-19
C58 VDD.n24 VSS 0.001388f
C59 VDD.n25 VSS 0.023172f
C60 VDD.t24 VSS 0.010883f
C61 VDD.t26 VSS 0.002466f
C62 VDD.n26 VSS 0.024709f
C63 VDD.t7 VSS 6.71e-19
C64 VDD.t3 VSS 6.71e-19
C65 VDD.n27 VSS 0.001388f
C66 VDD.n28 VSS 0.033097f
C67 VDD.t19 VSS 6.71e-19
C68 VDD.t13 VSS 6.71e-19
C69 VDD.n29 VSS 0.001388f
C70 VDD.n30 VSS 0.020255f
C71 VDD.t22 VSS 0.03828f
C72 VDD.t0 VSS 0.030576f
C73 VDD.t14 VSS 0.030576f
C74 VDD.t8 VSS 0.030576f
C75 VDD.t16 VSS 0.030576f
C76 VDD.t10 VSS 0.021984f
C77 VDD.t25 VSS 0.03828f
C78 VDD.t2 VSS 0.030576f
C79 VDD.t6 VSS 0.030576f
C80 VDD.t12 VSS 0.030576f
C81 VDD.t18 VSS 0.030576f
C82 VDD.t4 VSS 0.02388f
C83 VDD.n31 VSS -0.017931f
C84 VDD.t20 VSS 0.025145f
C85 VDD.n32 VSS 0.038891f
C86 VDD.n33 VSS 0.005278f
C87 VDD.t11 VSS 6.71e-19
C88 VDD.t5 VSS 6.71e-19
C89 VDD.n34 VSS 0.001388f
C90 VDD.n35 VSS 0.022776f
C91 VDD.n36 VSS 1.00176f
C92 INp.t4 VSS 0.192033f
C93 INp.t0 VSS 0.191404f
C94 INp.n0 VSS 0.237081f
C95 INp.t1 VSS 0.191404f
C96 INp.n1 VSS 0.139872f
C97 INp.t3 VSS 0.191404f
C98 INp.n2 VSS 0.121401f
C99 INp.t2 VSS 0.191893f
C100 INp.n3 VSS 0.332858f
C101 OUT.t11 VSS 0.007912f
C102 OUT.t9 VSS 0.007912f
C103 OUT.n0 VSS 0.018165f
C104 OUT.t10 VSS 0.007912f
C105 OUT.t2 VSS 0.007912f
C106 OUT.n1 VSS 0.023194f
C107 OUT.n2 VSS 0.320387f
C108 OUT.t7 VSS 0.007912f
C109 OUT.t5 VSS 0.007912f
C110 OUT.n3 VSS 0.018165f
C111 OUT.t1 VSS 0.007912f
C112 OUT.t4 VSS 0.007912f
C113 OUT.n4 VSS 0.023194f
C114 OUT.n5 VSS 0.306564f
C115 OUT.n6 VSS 0.848589f
C116 OUT.t8 VSS 0.007912f
C117 OUT.t6 VSS 0.007912f
C118 OUT.n7 VSS 0.018164f
C119 OUT.t0 VSS 0.007912f
C120 OUT.t3 VSS 0.007912f
C121 OUT.n8 VSS 0.023194f
C122 OUT.n9 VSS 0.303018f
C123 OUT.n10 VSS 0.376845f
.ends

