* NGSPICE file created from opamp_420.ext - technology: sky130A

.subckt opamp_nores OUT VSS VDD INp INn R
X0 a_320_185# VSS.t29 VSS.t30 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1 OUT.t10 INn.t0 a_578_185# VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2 VSS.t28 VSS.t26 VSS.t28 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X3 a_320_185# INp.t0 a_578_185# VSS.t5 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X4 VSS.t25 VSS.t22 VSS.t24 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0 ps=0 w=0.42 l=1
X5 a_320_185# a_320_185# VDD.t25 VDD.t24 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X6 a_578_185# R.t4 VSS.t8 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X7 VSS.t21 VSS.t20 OUT.t11 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X8 VSS.t3 R.t2 R.t3 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X9 VSS.t10 R.t5 a_578_185# VSS.t9 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X10 R.t1 R.t0 VSS.t34 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X11 VDD.t23 a_320_185# OUT.t3 VDD.t22 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X12 VDD.t21 a_320_185# a_320_185# VDD.t20 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X13 a_578_185# R.t6 VSS.t33 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X14 VDD.t19 a_320_185# OUT.t2 VDD.t18 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X15 OUT.t9 INn.t1 a_578_185# VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X16 a_320_185# VDD.t3 VDD.t5 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X17 OUT.t4 a_320_185# VDD.t17 VDD.t16 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X18 a_320_185# a_320_185# VDD.t15 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X19 a_578_185# INp.t1 a_320_185# VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X20 VDD.t2 VDD.t0 OUT.t5 VDD.t1 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X21 a_578_185# INp.t2 a_320_185# VSS.t27 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X22 OUT.t8 INn.t2 a_578_185# VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X23 VSS.t19 VSS.t17 VSS.t19 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X24 VSS.t16 VSS.t15 VSS.t16 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X25 VSS.t31 R.t7 a_578_185# VSS.t5 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X26 VSS.t14 VSS.t13 VSS.t14 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X27 a_320_185# INp.t3 a_578_185# VSS.t9 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X28 OUT.t0 a_320_185# VDD.t13 VDD.t12 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X29 a_578_185# INn.t3 OUT.t7 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X30 a_578_185# INp.t4 a_320_185# VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X31 VDD.t11 a_320_185# a_320_185# VDD.t10 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X32 a_578_185# INn.t4 OUT.t6 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X33 VDD.t9 a_320_185# a_320_185# VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X34 OUT.t1 a_320_185# VDD.t7 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X35 VSS.t12 VSS.t11 VSS.t12 VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
R0 VSS.t23 VSS.t18 128418
R1 VSS.t18 VSS.t0 1051.11
R2 VSS.t0 VSS.t4 1051.11
R3 VSS.t4 VSS.t5 1051.11
R4 VSS.t5 VSS.t7 1051.11
R5 VSS.t7 VSS.t2 1051.11
R6 VSS.t6 VSS.t9 1051.11
R7 VSS.t9 VSS.t32 1051.11
R8 VSS.t32 VSS.t1 1051.11
R9 VSS.t1 VSS.t27 1051.11
R10 VSS.t27 VSS.t23 1051.11
R11 VSS.n26 VSS.t2 541.852
R12 VSS.n26 VSS.t6 509.26
R13 VSS.t19 VSS.n3 235.764
R14 VSS.n15 VSS.t25 235.763
R15 VSS.n23 VSS.n22 194.573
R16 VSS.n10 VSS.n9 194.542
R17 VSS.n25 VSS.n24 194.463
R18 VSS.n12 VSS.n11 194.463
R19 VSS.n18 VSS.n17 194.3
R20 VSS.n21 VSS.n20 194.3
R21 VSS.n8 VSS.n7 194.3
R22 VSS.n5 VSS.n4 194.3
R23 VSS.n14 VSS.t29 118.005
R24 VSS.n2 VSS.t20 118.005
R25 VSS.n16 VSS.t22 104.028
R26 VSS.n19 VSS.t26 104.028
R27 VSS.n13 VSS.t11 104.028
R28 VSS.n0 VSS.t13 104.028
R29 VSS.n6 VSS.t15 104.028
R30 VSS.n1 VSS.t17 104.028
R31 VSS.n14 VSS.t30 87.6949
R32 VSS.n2 VSS.t21 87.5315
R33 VSS.n22 VSS.t33 41.4291
R34 VSS.n22 VSS.t12 41.4291
R35 VSS.n17 VSS.t28 41.4291
R36 VSS.n17 VSS.t24 41.4291
R37 VSS.t12 VSS.n21 41.4291
R38 VSS.n21 VSS.t28 41.4291
R39 VSS.n24 VSS.t34 41.4291
R40 VSS.n24 VSS.t10 41.4291
R41 VSS.n9 VSS.t14 41.4291
R42 VSS.n9 VSS.t31 41.4291
R43 VSS.n8 VSS.t16 41.4291
R44 VSS.t14 VSS.n8 41.4291
R45 VSS.n4 VSS.t19 41.4291
R46 VSS.n4 VSS.t16 41.4291
R47 VSS.n11 VSS.t8 41.4291
R48 VSS.n11 VSS.t3 41.4291
R49 VSS.n27 VSS.n26 26.2219
R50 VSS.n25 VSS.n23 0.728909
R51 VSS.n12 VSS.n10 0.690273
R52 VSS VSS.n28 0.314125
R53 VSS.n28 VSS.n12 0.216409
R54 VSS.n27 VSS.n25 0.210727
R55 VSS.n20 VSS.n13 0.0429342
R56 VSS.n20 VSS.n19 0.0429342
R57 VSS.n19 VSS.n18 0.0429342
R58 VSS.n18 VSS.n16 0.0429342
R59 VSS.n5 VSS.n1 0.0429342
R60 VSS.n6 VSS.n5 0.0429342
R61 VSS.n7 VSS.n6 0.0429342
R62 VSS.n7 VSS.n0 0.0429342
R63 VSS.n15 VSS.n14 0.0405
R64 VSS.n3 VSS.n2 0.0389615
R65 VSS.n23 VSS.n13 0.0347105
R66 VSS.n10 VSS.n0 0.0340526
R67 VSS.n16 VSS.n15 0.00872368
R68 VSS.n3 VSS.n1 0.00773684
R69 VSS.n28 VSS.n27 0.00618182
R70 INn.n0 INn.t1 118.769
R71 INn.n3 INn.t2 118.005
R72 INn.n2 INn.t3 118.005
R73 INn.n1 INn.t0 118.005
R74 INn.n0 INn.t4 118.005
R75 INn INn.n3 3.33334
R76 INn.n1 INn.n0 2.66195
R77 INn.n3 INn.n2 2.55325
R78 INn.n2 INn.n1 0.764886
R79 OUT.n9 OUT.n7 204.206
R80 OUT.n5 OUT.n3 204.206
R81 OUT.n2 OUT.n0 204.206
R82 OUT.n9 OUT.n8 71.1729
R83 OUT.n5 OUT.n4 71.1729
R84 OUT.n2 OUT.n1 71.1729
R85 OUT.n7 OUT.t2 28.5655
R86 OUT.n7 OUT.t0 28.5655
R87 OUT.n3 OUT.t3 28.5655
R88 OUT.n3 OUT.t4 28.5655
R89 OUT.n0 OUT.t5 28.5655
R90 OUT.n0 OUT.t1 28.5655
R91 OUT.n8 OUT.t6 17.4005
R92 OUT.n8 OUT.t9 17.4005
R93 OUT.n4 OUT.t7 17.4005
R94 OUT.n4 OUT.t10 17.4005
R95 OUT.n1 OUT.t11 17.4005
R96 OUT.n1 OUT.t8 17.4005
R97 OUT.n6 OUT.n2 3.7629
R98 OUT.n6 OUT.n5 3.4105
R99 OUT.n10 OUT.n9 3.4105
R100 OUT.n10 OUT.n6 0.19414
R101 OUT OUT.n10 0.0146
R102 INp.n0 INp.t4 118.769
R103 INp.n3 INp.t2 118.621
R104 INp.n2 INp.t3 118.005
R105 INp.n1 INp.t1 118.005
R106 INp.n0 INp.t0 118.005
R107 INp INp.n3 2.77717
R108 INp.n1 INp.n0 2.66195
R109 INp.n3 INp.n2 1.71868
R110 INp.n2 INp.n1 0.764886
R111 VDD.t6 VDD.t1 478.712
R112 VDD.t20 VDD.t6 478.712
R113 VDD.t14 VDD.t20 478.712
R114 VDD.t22 VDD.t14 478.712
R115 VDD.t16 VDD.t22 478.712
R116 VDD.t10 VDD.t24 478.712
R117 VDD.t24 VDD.t18 478.712
R118 VDD.t18 VDD.t12 478.712
R119 VDD.t12 VDD.t8 478.712
R120 VDD.t8 VDD.t4 478.712
R121 VDD.n10 VDD.t10 269.043
R122 VDD.n5 VDD.t5 228.215
R123 VDD.n0 VDD.t2 228.215
R124 VDD.n10 VDD.t16 209.668
R125 VDD.n7 VDD.n6 199.851
R126 VDD.n9 VDD.n8 199.851
R127 VDD.n2 VDD.n1 199.851
R128 VDD.n4 VDD.n3 199.851
R129 VDD.n13 VDD.n12 199.851
R130 VDD.n0 VDD.t0 120.855
R131 VDD.n5 VDD.t3 120.749
R132 VDD.n11 VDD.n10 38.9956
R133 VDD.n6 VDD.t13 28.5655
R134 VDD.n6 VDD.t9 28.5655
R135 VDD.n8 VDD.t25 28.5655
R136 VDD.n8 VDD.t19 28.5655
R137 VDD.n1 VDD.t7 28.5655
R138 VDD.n1 VDD.t21 28.5655
R139 VDD.n3 VDD.t15 28.5655
R140 VDD.n3 VDD.t23 28.5655
R141 VDD.n12 VDD.t17 28.5655
R142 VDD.n12 VDD.t11 28.5655
R143 VDD.n2 VDD.n0 0.890989
R144 VDD.n7 VDD.n5 0.760446
R145 VDD.n9 VDD.n7 0.40675
R146 VDD.n4 VDD.n2 0.40675
R147 VDD.n13 VDD.n4 0.40675
R148 VDD VDD.n13 0.357528
R149 VDD.n13 VDD.n11 0.208833
R150 VDD.n11 VDD.n9 0.188
R151 R.n5 R.n0 194.387
R152 R.n3 R.t6 104.575
R153 R.n1 R.t7 104.575
R154 R.n3 R.t5 104.028
R155 R.n4 R.t0 104.028
R156 R.n2 R.t2 104.028
R157 R.n1 R.t4 104.028
R158 R.n0 R.t3 41.4291
R159 R.n0 R.t1 41.4291
R160 R R.n5 3.54374
R161 R.n4 R.n3 0.54711
R162 R.n2 R.n1 0.54711
R163 R.n5 R.n4 0.171686
R164 R.n5 R.n2 0.167449
.ends

