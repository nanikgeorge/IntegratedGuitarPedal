magic
tech sky130A
magscale 1 2
timestamp 1713395545
<< pwell >>
rect -425 -279 425 279
<< nmos >>
rect -229 -69 -29 131
rect 29 -69 229 131
<< ndiff >>
rect -287 119 -229 131
rect -287 -57 -275 119
rect -241 -57 -229 119
rect -287 -69 -229 -57
rect -29 119 29 131
rect -29 -57 -17 119
rect 17 -57 29 119
rect -29 -69 29 -57
rect 229 119 287 131
rect 229 -57 241 119
rect 275 -57 287 119
rect 229 -69 287 -57
<< ndiffc >>
rect -275 -57 -241 119
rect -17 -57 17 119
rect 241 -57 275 119
<< psubdiff >>
rect -389 209 389 243
rect -389 147 -355 209
rect 355 147 389 209
rect -389 -209 -355 -147
rect 355 -209 389 -147
rect -389 -243 -293 -209
rect 293 -243 389 -209
<< psubdiffcont >>
rect -389 -147 -355 147
rect 355 -147 389 147
rect -293 -243 293 -209
<< poly >>
rect -229 131 -29 157
rect 29 131 229 157
rect -229 -107 -29 -69
rect -229 -141 -213 -107
rect -45 -141 -29 -107
rect -229 -157 -29 -141
rect 29 -107 229 -69
rect 29 -141 45 -107
rect 213 -141 229 -107
rect 29 -157 229 -141
<< polycont >>
rect -213 -141 -45 -107
rect 45 -141 213 -107
<< locali >>
rect -389 147 -355 163
rect 355 147 389 163
rect -275 119 -241 135
rect -275 -73 -241 -57
rect -17 119 17 135
rect -17 -73 17 -57
rect 241 119 275 135
rect 241 -73 275 -57
rect -229 -141 -213 -107
rect -45 -141 -29 -107
rect 29 -141 45 -107
rect 213 -141 229 -107
rect -389 -163 -355 -147
rect 355 -163 389 -147
rect -309 -243 -293 -209
rect 293 -243 309 -209
<< viali >>
rect -275 -57 -241 119
rect -17 -57 17 119
rect 241 -57 275 119
rect -213 -141 -45 -107
rect 45 -141 213 -107
<< metal1 >>
rect -281 119 -235 131
rect -281 -57 -275 119
rect -241 -57 -235 119
rect -281 -69 -235 -57
rect -23 119 23 131
rect -23 -57 -17 119
rect 17 -57 23 119
rect -23 -69 23 -57
rect 235 119 281 131
rect 235 -57 241 119
rect 275 -57 281 119
rect 235 -69 281 -57
rect -225 -107 -33 -101
rect -225 -141 -213 -107
rect -45 -141 -33 -107
rect -225 -147 -33 -141
rect 33 -107 225 -101
rect 33 -141 45 -107
rect 213 -141 225 -107
rect 33 -147 225 -141
<< properties >>
string FIXED_BBOX -372 -226 372 226
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 1 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
