MACRO tt_um_guitar_pedal
  CLASS BLOCK ;
  FOREIGN tt_um_guitar_pedal ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.000000 ;
    ANTENNADIFFAREA 0.870000 ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.740000 ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 5.000 5.000 6.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 157.530 5.000 159.030 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 27.950 188.800 56.450 189.800 ;
        RECT 27.950 176.800 28.950 188.800 ;
      LAYER pwell ;
        RECT 29.450 187.300 54.950 188.300 ;
        RECT 29.450 178.300 36.900 187.300 ;
      LAYER nwell ;
        RECT 37.080 183.860 53.210 186.420 ;
      LAYER pwell ;
        RECT 37.050 179.450 53.200 180.300 ;
        RECT 53.950 178.300 54.950 187.300 ;
        RECT 29.450 177.300 54.950 178.300 ;
      LAYER nwell ;
        RECT 55.450 176.800 56.450 188.800 ;
        RECT 63.485 189.625 67.735 192.465 ;
        RECT 27.950 175.800 56.450 176.800 ;
      LAYER pwell ;
        RECT 47.150 172.900 56.970 174.910 ;
        RECT 57.350 172.900 59.360 188.720 ;
        RECT 63.485 186.835 67.735 189.625 ;
      LAYER nwell ;
        RECT 92.020 189.580 120.520 190.580 ;
        RECT 63.485 182.325 67.735 185.165 ;
      LAYER pwell ;
        RECT 63.485 179.535 67.735 182.325 ;
      LAYER nwell ;
        RECT 92.020 177.580 93.020 189.580 ;
      LAYER pwell ;
        RECT 93.520 188.080 119.020 189.080 ;
        RECT 93.520 179.080 100.970 188.080 ;
      LAYER nwell ;
        RECT 101.150 184.640 117.280 187.200 ;
      LAYER pwell ;
        RECT 101.120 180.230 117.270 181.080 ;
        RECT 118.020 179.080 119.020 188.080 ;
        RECT 93.520 178.080 119.020 179.080 ;
      LAYER nwell ;
        RECT 119.520 177.580 120.520 189.580 ;
        RECT 127.555 190.405 131.805 193.245 ;
        RECT 62.450 175.645 67.890 177.250 ;
        RECT 92.020 176.580 120.520 177.580 ;
      LAYER pwell ;
        RECT 62.810 174.445 66.680 175.355 ;
        RECT 66.795 174.530 67.685 175.315 ;
        RECT 62.810 174.425 62.955 174.445 ;
        RECT 62.785 174.255 62.955 174.425 ;
        RECT 111.220 173.680 121.040 175.690 ;
        RECT 121.420 173.680 123.430 189.500 ;
        RECT 127.555 187.615 131.805 190.405 ;
      LAYER nwell ;
        RECT 127.555 183.105 131.805 185.945 ;
      LAYER pwell ;
        RECT 127.555 180.315 131.805 183.105 ;
      LAYER nwell ;
        RECT 126.520 176.425 131.960 178.030 ;
      LAYER pwell ;
        RECT 126.880 175.225 130.750 176.135 ;
        RECT 130.865 175.310 131.755 176.095 ;
        RECT 126.880 175.205 127.025 175.225 ;
        RECT 126.855 175.035 127.025 175.205 ;
      LAYER nwell ;
        RECT 28.180 159.360 56.680 160.360 ;
        RECT 28.180 147.360 29.180 159.360 ;
      LAYER pwell ;
        RECT 29.680 157.860 55.180 158.860 ;
        RECT 29.680 148.860 37.130 157.860 ;
      LAYER nwell ;
        RECT 37.310 154.420 53.440 156.980 ;
      LAYER pwell ;
        RECT 37.280 150.010 53.430 150.860 ;
        RECT 54.180 148.860 55.180 157.860 ;
        RECT 29.680 147.860 55.180 148.860 ;
      LAYER nwell ;
        RECT 55.680 147.360 56.680 159.360 ;
        RECT 63.715 160.185 67.965 163.025 ;
        RECT 28.180 146.360 56.680 147.360 ;
      LAYER pwell ;
        RECT 47.380 143.460 57.200 145.470 ;
        RECT 57.580 143.460 59.590 159.280 ;
        RECT 63.715 157.395 67.965 160.185 ;
      LAYER nwell ;
        RECT 91.840 158.980 120.340 159.980 ;
        RECT 63.715 152.885 67.965 155.725 ;
      LAYER pwell ;
        RECT 63.715 150.095 67.965 152.885 ;
      LAYER nwell ;
        RECT 62.680 146.205 68.120 147.810 ;
        RECT 91.840 146.980 92.840 158.980 ;
      LAYER pwell ;
        RECT 93.340 157.480 118.840 158.480 ;
        RECT 93.340 148.480 100.790 157.480 ;
      LAYER nwell ;
        RECT 100.970 154.040 117.100 156.600 ;
      LAYER pwell ;
        RECT 100.940 149.630 117.090 150.480 ;
        RECT 117.840 148.480 118.840 157.480 ;
        RECT 93.340 147.480 118.840 148.480 ;
      LAYER nwell ;
        RECT 119.340 146.980 120.340 158.980 ;
        RECT 127.375 159.805 131.625 162.645 ;
        RECT 91.840 145.980 120.340 146.980 ;
      LAYER pwell ;
        RECT 63.040 145.005 66.910 145.915 ;
        RECT 67.025 145.090 67.915 145.875 ;
        RECT 63.040 144.985 63.185 145.005 ;
        RECT 63.015 144.815 63.185 144.985 ;
        RECT 111.040 143.080 120.860 145.090 ;
        RECT 121.240 143.080 123.250 158.900 ;
        RECT 127.375 157.015 131.625 159.805 ;
      LAYER nwell ;
        RECT 127.375 152.505 131.625 155.345 ;
      LAYER pwell ;
        RECT 127.375 149.715 131.625 152.505 ;
      LAYER nwell ;
        RECT 126.340 145.825 131.780 147.430 ;
      LAYER pwell ;
        RECT 126.700 144.625 130.570 145.535 ;
        RECT 130.685 144.710 131.575 145.495 ;
        RECT 126.700 144.605 126.845 144.625 ;
        RECT 126.675 144.435 126.845 144.605 ;
      LAYER nwell ;
        RECT 28.780 125.840 57.280 126.840 ;
        RECT 28.780 113.840 29.780 125.840 ;
      LAYER pwell ;
        RECT 30.280 124.340 55.780 125.340 ;
        RECT 30.280 115.340 37.730 124.340 ;
      LAYER nwell ;
        RECT 37.910 120.900 54.040 123.460 ;
      LAYER pwell ;
        RECT 37.880 116.490 54.030 117.340 ;
        RECT 54.780 115.340 55.780 124.340 ;
        RECT 30.280 114.340 55.780 115.340 ;
      LAYER nwell ;
        RECT 56.280 113.840 57.280 125.840 ;
        RECT 64.315 126.665 68.565 129.505 ;
        RECT 28.780 112.840 57.280 113.840 ;
      LAYER pwell ;
        RECT 47.980 109.940 57.800 111.950 ;
        RECT 58.180 109.940 60.190 125.760 ;
        RECT 64.315 123.875 68.565 126.665 ;
      LAYER nwell ;
        RECT 92.320 125.190 120.820 126.190 ;
        RECT 64.315 119.365 68.565 122.205 ;
      LAYER pwell ;
        RECT 64.315 116.575 68.565 119.365 ;
      LAYER nwell ;
        RECT 63.280 112.685 68.720 114.290 ;
        RECT 92.320 113.190 93.320 125.190 ;
      LAYER pwell ;
        RECT 93.820 123.690 119.320 124.690 ;
        RECT 93.820 114.690 101.270 123.690 ;
      LAYER nwell ;
        RECT 101.450 120.250 117.580 122.810 ;
      LAYER pwell ;
        RECT 101.420 115.840 117.570 116.690 ;
        RECT 118.320 114.690 119.320 123.690 ;
        RECT 93.820 113.690 119.320 114.690 ;
      LAYER nwell ;
        RECT 119.820 113.190 120.820 125.190 ;
        RECT 127.855 126.015 132.105 128.855 ;
      LAYER pwell ;
        RECT 63.640 111.485 67.510 112.395 ;
        RECT 67.625 111.570 68.515 112.355 ;
      LAYER nwell ;
        RECT 92.320 112.190 120.820 113.190 ;
      LAYER pwell ;
        RECT 63.640 111.465 63.785 111.485 ;
        RECT 63.615 111.295 63.785 111.465 ;
        RECT 111.520 109.290 121.340 111.300 ;
        RECT 121.720 109.290 123.730 125.110 ;
        RECT 127.855 123.225 132.105 126.015 ;
      LAYER nwell ;
        RECT 127.855 118.715 132.105 121.555 ;
      LAYER pwell ;
        RECT 127.855 115.925 132.105 118.715 ;
      LAYER nwell ;
        RECT 126.820 112.035 132.260 113.640 ;
      LAYER pwell ;
        RECT 127.180 110.835 131.050 111.745 ;
        RECT 131.165 110.920 132.055 111.705 ;
        RECT 127.180 110.815 127.325 110.835 ;
        RECT 127.155 110.645 127.325 110.815 ;
      LAYER nwell ;
        RECT 28.160 90.610 56.660 91.610 ;
        RECT 28.160 78.610 29.160 90.610 ;
      LAYER pwell ;
        RECT 29.660 89.110 55.160 90.110 ;
        RECT 29.660 80.110 37.110 89.110 ;
      LAYER nwell ;
        RECT 37.290 85.670 53.420 88.230 ;
      LAYER pwell ;
        RECT 37.260 81.260 53.410 82.110 ;
        RECT 54.160 80.110 55.160 89.110 ;
        RECT 29.660 79.110 55.160 80.110 ;
      LAYER nwell ;
        RECT 55.660 78.610 56.660 90.610 ;
        RECT 63.695 91.435 67.945 94.275 ;
        RECT 28.160 77.610 56.660 78.610 ;
      LAYER pwell ;
        RECT 47.360 74.710 57.180 76.720 ;
        RECT 57.560 74.710 59.570 90.530 ;
        RECT 63.695 88.645 67.945 91.435 ;
      LAYER nwell ;
        RECT 94.070 89.960 122.570 90.960 ;
        RECT 63.695 84.135 67.945 86.975 ;
      LAYER pwell ;
        RECT 63.695 81.345 67.945 84.135 ;
      LAYER nwell ;
        RECT 62.660 77.455 68.100 79.060 ;
        RECT 94.070 77.960 95.070 89.960 ;
      LAYER pwell ;
        RECT 95.570 88.460 121.070 89.460 ;
        RECT 95.570 79.460 103.020 88.460 ;
      LAYER nwell ;
        RECT 103.200 85.020 119.330 87.580 ;
      LAYER pwell ;
        RECT 103.170 80.610 119.320 81.460 ;
        RECT 120.070 79.460 121.070 88.460 ;
        RECT 95.570 78.460 121.070 79.460 ;
      LAYER nwell ;
        RECT 121.570 77.960 122.570 89.960 ;
        RECT 129.605 90.785 133.855 93.625 ;
      LAYER pwell ;
        RECT 63.020 76.255 66.890 77.165 ;
        RECT 67.005 76.340 67.895 77.125 ;
      LAYER nwell ;
        RECT 94.070 76.960 122.570 77.960 ;
      LAYER pwell ;
        RECT 63.020 76.235 63.165 76.255 ;
        RECT 62.995 76.065 63.165 76.235 ;
        RECT 113.270 74.060 123.090 76.070 ;
        RECT 123.470 74.060 125.480 89.880 ;
        RECT 129.605 87.995 133.855 90.785 ;
      LAYER nwell ;
        RECT 129.605 83.485 133.855 86.325 ;
      LAYER pwell ;
        RECT 129.605 80.695 133.855 83.485 ;
      LAYER nwell ;
        RECT 128.570 76.805 134.010 78.410 ;
      LAYER pwell ;
        RECT 128.930 75.605 132.800 76.515 ;
        RECT 132.915 75.690 133.805 76.475 ;
        RECT 128.930 75.585 129.075 75.605 ;
        RECT 128.905 75.415 129.075 75.585 ;
      LAYER li1 ;
        RECT 127.570 192.880 131.820 193.130 ;
        RECT 63.500 192.100 67.750 192.350 ;
        RECT 63.500 190.100 63.850 192.100 ;
        RECT 64.465 191.600 65.465 191.770 ;
        RECT 65.755 191.600 66.755 191.770 ;
        RECT 67.350 191.500 67.750 192.100 ;
        RECT 64.235 191.350 64.405 191.385 ;
        RECT 64.150 190.500 64.500 191.350 ;
        RECT 64.150 190.100 65.150 190.500 ;
        RECT 65.525 190.345 65.695 191.385 ;
        RECT 66.815 191.350 66.985 191.385 ;
        RECT 66.750 190.500 67.050 191.350 ;
        RECT 64.850 189.700 65.150 190.100 ;
        RECT 66.050 190.100 67.050 190.500 ;
        RECT 67.350 190.200 68.750 191.500 ;
        RECT 127.570 190.880 127.920 192.880 ;
        RECT 128.535 192.380 129.535 192.550 ;
        RECT 129.825 192.380 130.825 192.550 ;
        RECT 131.420 192.280 131.820 192.880 ;
        RECT 128.305 192.130 128.475 192.165 ;
        RECT 128.220 191.280 128.570 192.130 ;
        RECT 128.220 190.880 129.220 191.280 ;
        RECT 129.595 191.125 129.765 192.165 ;
        RECT 130.885 192.130 131.055 192.165 ;
        RECT 130.820 191.280 131.120 192.130 ;
        RECT 128.920 190.480 129.220 190.880 ;
        RECT 130.120 190.880 131.120 191.280 ;
        RECT 131.420 190.980 132.820 192.280 ;
        RECT 130.120 190.480 130.420 190.880 ;
        RECT 66.050 189.700 66.350 190.100 ;
        RECT 28.370 189.220 56.090 189.550 ;
        RECT 64.850 189.300 66.350 189.700 ;
        RECT 92.440 190.000 120.160 190.330 ;
        RECT 128.920 190.080 130.420 190.480 ;
        RECT 28.370 176.350 28.700 189.220 ;
        RECT 29.690 187.570 54.770 187.900 ;
        RECT 29.690 178.000 30.020 187.570 ;
        RECT 34.550 185.600 53.000 186.200 ;
        RECT 37.320 184.340 37.490 185.380 ;
        RECT 38.610 184.340 38.780 185.380 ;
        RECT 39.900 184.340 40.070 185.380 ;
        RECT 41.190 184.340 41.360 185.380 ;
        RECT 42.480 184.340 42.650 185.380 ;
        RECT 43.770 184.340 43.940 185.380 ;
        RECT 45.060 184.340 45.230 185.380 ;
        RECT 46.350 184.340 46.520 185.380 ;
        RECT 47.640 184.340 47.810 185.380 ;
        RECT 48.930 184.340 49.100 185.380 ;
        RECT 50.220 184.340 50.390 185.380 ;
        RECT 51.510 184.340 51.680 185.380 ;
        RECT 52.800 184.340 52.970 185.380 ;
        RECT 37.550 183.955 38.550 184.125 ;
        RECT 38.840 183.955 39.840 184.125 ;
        RECT 40.130 183.955 41.130 184.125 ;
        RECT 41.420 183.955 42.420 184.125 ;
        RECT 42.710 183.955 43.710 184.125 ;
        RECT 44.000 183.955 45.000 184.125 ;
        RECT 45.290 183.955 46.290 184.125 ;
        RECT 46.580 183.955 47.580 184.125 ;
        RECT 47.870 183.955 48.870 184.125 ;
        RECT 49.160 183.955 50.160 184.125 ;
        RECT 50.450 183.955 51.450 184.125 ;
        RECT 51.740 183.955 52.740 184.125 ;
        RECT 38.840 183.415 39.840 183.585 ;
        RECT 42.710 183.415 43.710 183.585 ;
        RECT 44.000 183.415 45.000 183.585 ;
        RECT 47.870 183.415 48.870 183.585 ;
        RECT 49.160 183.415 50.160 183.585 ;
        RECT 37.320 182.205 37.490 183.245 ;
        RECT 38.610 182.205 38.780 183.245 ;
        RECT 39.900 182.205 40.070 183.245 ;
        RECT 41.190 182.205 41.360 183.245 ;
        RECT 42.480 182.205 42.650 183.245 ;
        RECT 43.770 182.205 43.940 183.245 ;
        RECT 45.060 182.205 45.230 183.245 ;
        RECT 46.350 182.205 46.520 183.245 ;
        RECT 47.640 182.205 47.810 183.245 ;
        RECT 48.930 182.205 49.100 183.245 ;
        RECT 50.220 182.205 50.390 183.245 ;
        RECT 51.510 182.205 51.680 183.245 ;
        RECT 52.800 182.205 52.970 183.245 ;
        RECT 37.550 181.865 38.550 182.035 ;
        RECT 40.130 181.865 41.130 182.035 ;
        RECT 41.420 181.865 42.420 182.035 ;
        RECT 45.290 181.865 46.290 182.035 ;
        RECT 46.580 181.865 47.580 182.035 ;
        RECT 50.450 181.865 51.450 182.035 ;
        RECT 51.740 181.865 52.740 182.035 ;
        RECT 37.550 181.235 38.550 181.405 ;
        RECT 38.840 181.235 39.840 181.405 ;
        RECT 40.130 181.235 41.130 181.405 ;
        RECT 41.420 181.235 42.420 181.405 ;
        RECT 42.710 181.235 43.710 181.405 ;
        RECT 44.000 181.235 45.000 181.405 ;
        RECT 45.290 181.235 46.290 181.405 ;
        RECT 46.580 181.235 47.580 181.405 ;
        RECT 47.870 181.235 48.870 181.405 ;
        RECT 49.160 181.235 50.160 181.405 ;
        RECT 50.450 181.235 51.450 181.405 ;
        RECT 51.740 181.235 52.740 181.405 ;
        RECT 37.320 180.605 37.490 181.065 ;
        RECT 38.610 180.605 38.780 181.065 ;
        RECT 39.900 180.605 40.070 181.065 ;
        RECT 41.190 180.605 41.360 181.065 ;
        RECT 42.480 180.605 42.650 181.065 ;
        RECT 43.770 180.605 43.940 181.065 ;
        RECT 45.060 180.605 45.230 181.065 ;
        RECT 46.350 180.605 46.520 181.065 ;
        RECT 47.640 180.605 47.810 181.065 ;
        RECT 48.930 180.605 49.100 181.065 ;
        RECT 50.220 180.605 50.390 181.065 ;
        RECT 51.510 180.605 51.680 181.065 ;
        RECT 52.800 180.605 52.970 181.065 ;
        RECT 34.550 179.800 36.750 180.500 ;
        RECT 37.300 179.650 53.000 180.200 ;
        RECT 54.440 178.000 54.770 187.570 ;
        RECT 29.690 177.670 54.770 178.000 ;
        RECT 55.760 176.350 56.090 189.220 ;
        RECT 57.530 188.370 59.180 188.540 ;
        RECT 57.530 180.200 57.700 188.370 ;
        RECT 57.950 185.700 58.750 187.900 ;
        RECT 56.950 177.800 57.700 180.200 ;
        RECT 28.370 176.020 56.090 176.350 ;
        RECT 47.450 174.730 53.250 175.200 ;
        RECT 47.330 174.700 56.790 174.730 ;
        RECT 57.530 174.700 57.700 177.800 ;
        RECT 47.330 174.560 57.700 174.700 ;
        RECT 47.330 173.250 47.500 174.560 ;
        RECT 47.980 173.730 50.140 174.080 ;
        RECT 53.980 173.730 56.140 174.080 ;
        RECT 56.620 173.250 57.700 174.560 ;
        RECT 58.180 173.730 58.530 175.890 ;
        RECT 59.010 173.250 59.180 188.370 ;
        RECT 63.500 187.200 63.850 189.100 ;
        RECT 64.150 188.100 64.500 189.100 ;
        RECT 64.235 187.865 64.405 188.100 ;
        RECT 65.350 187.900 65.850 189.300 ;
        RECT 66.750 188.100 67.050 189.100 ;
        RECT 65.525 187.865 65.695 187.900 ;
        RECT 66.815 187.865 66.985 188.100 ;
        RECT 67.350 187.800 68.750 189.100 ;
        RECT 64.465 187.525 65.465 187.695 ;
        RECT 65.755 187.525 66.755 187.695 ;
        RECT 67.350 187.200 67.750 187.800 ;
        RECT 63.500 186.850 67.750 187.200 ;
        RECT 63.500 184.800 67.750 185.050 ;
        RECT 63.500 182.800 63.850 184.800 ;
        RECT 64.465 184.300 65.465 184.470 ;
        RECT 65.755 184.300 66.755 184.470 ;
        RECT 67.350 184.200 67.750 184.800 ;
        RECT 64.235 184.050 64.405 184.085 ;
        RECT 64.150 183.200 64.500 184.050 ;
        RECT 64.150 182.800 65.150 183.200 ;
        RECT 65.525 183.045 65.695 184.085 ;
        RECT 66.815 184.050 66.985 184.085 ;
        RECT 66.750 183.200 67.050 184.050 ;
        RECT 64.850 182.400 65.150 182.800 ;
        RECT 66.050 182.800 67.050 183.200 ;
        RECT 67.350 182.900 68.750 184.200 ;
        RECT 66.050 182.400 66.350 182.800 ;
        RECT 64.850 182.000 66.350 182.400 ;
        RECT 63.500 179.900 63.850 181.800 ;
        RECT 64.150 180.800 64.500 181.800 ;
        RECT 64.235 180.565 64.405 180.800 ;
        RECT 65.350 180.600 65.850 182.000 ;
        RECT 66.750 180.800 67.050 181.800 ;
        RECT 65.525 180.565 65.695 180.600 ;
        RECT 66.815 180.565 66.985 180.800 ;
        RECT 67.350 180.500 68.750 181.800 ;
        RECT 64.465 180.225 65.465 180.395 ;
        RECT 65.755 180.225 66.755 180.395 ;
        RECT 67.350 179.900 67.750 180.500 ;
        RECT 63.500 179.550 67.750 179.900 ;
        RECT 62.640 176.975 67.700 177.145 ;
        RECT 92.440 177.130 92.770 190.000 ;
        RECT 93.760 188.350 118.840 188.680 ;
        RECT 93.760 178.780 94.090 188.350 ;
        RECT 98.620 186.380 117.070 186.980 ;
        RECT 101.390 185.120 101.560 186.160 ;
        RECT 102.680 185.120 102.850 186.160 ;
        RECT 103.970 185.120 104.140 186.160 ;
        RECT 105.260 185.120 105.430 186.160 ;
        RECT 106.550 185.120 106.720 186.160 ;
        RECT 107.840 185.120 108.010 186.160 ;
        RECT 109.130 185.120 109.300 186.160 ;
        RECT 110.420 185.120 110.590 186.160 ;
        RECT 111.710 185.120 111.880 186.160 ;
        RECT 113.000 185.120 113.170 186.160 ;
        RECT 114.290 185.120 114.460 186.160 ;
        RECT 115.580 185.120 115.750 186.160 ;
        RECT 116.870 185.120 117.040 186.160 ;
        RECT 101.620 184.735 102.620 184.905 ;
        RECT 102.910 184.735 103.910 184.905 ;
        RECT 104.200 184.735 105.200 184.905 ;
        RECT 105.490 184.735 106.490 184.905 ;
        RECT 106.780 184.735 107.780 184.905 ;
        RECT 108.070 184.735 109.070 184.905 ;
        RECT 109.360 184.735 110.360 184.905 ;
        RECT 110.650 184.735 111.650 184.905 ;
        RECT 111.940 184.735 112.940 184.905 ;
        RECT 113.230 184.735 114.230 184.905 ;
        RECT 114.520 184.735 115.520 184.905 ;
        RECT 115.810 184.735 116.810 184.905 ;
        RECT 102.910 184.195 103.910 184.365 ;
        RECT 106.780 184.195 107.780 184.365 ;
        RECT 108.070 184.195 109.070 184.365 ;
        RECT 111.940 184.195 112.940 184.365 ;
        RECT 113.230 184.195 114.230 184.365 ;
        RECT 101.390 182.985 101.560 184.025 ;
        RECT 102.680 182.985 102.850 184.025 ;
        RECT 103.970 182.985 104.140 184.025 ;
        RECT 105.260 182.985 105.430 184.025 ;
        RECT 106.550 182.985 106.720 184.025 ;
        RECT 107.840 182.985 108.010 184.025 ;
        RECT 109.130 182.985 109.300 184.025 ;
        RECT 110.420 182.985 110.590 184.025 ;
        RECT 111.710 182.985 111.880 184.025 ;
        RECT 113.000 182.985 113.170 184.025 ;
        RECT 114.290 182.985 114.460 184.025 ;
        RECT 115.580 182.985 115.750 184.025 ;
        RECT 116.870 182.985 117.040 184.025 ;
        RECT 101.620 182.645 102.620 182.815 ;
        RECT 104.200 182.645 105.200 182.815 ;
        RECT 105.490 182.645 106.490 182.815 ;
        RECT 109.360 182.645 110.360 182.815 ;
        RECT 110.650 182.645 111.650 182.815 ;
        RECT 114.520 182.645 115.520 182.815 ;
        RECT 115.810 182.645 116.810 182.815 ;
        RECT 101.620 182.015 102.620 182.185 ;
        RECT 102.910 182.015 103.910 182.185 ;
        RECT 104.200 182.015 105.200 182.185 ;
        RECT 105.490 182.015 106.490 182.185 ;
        RECT 106.780 182.015 107.780 182.185 ;
        RECT 108.070 182.015 109.070 182.185 ;
        RECT 109.360 182.015 110.360 182.185 ;
        RECT 110.650 182.015 111.650 182.185 ;
        RECT 111.940 182.015 112.940 182.185 ;
        RECT 113.230 182.015 114.230 182.185 ;
        RECT 114.520 182.015 115.520 182.185 ;
        RECT 115.810 182.015 116.810 182.185 ;
        RECT 101.390 181.385 101.560 181.845 ;
        RECT 102.680 181.385 102.850 181.845 ;
        RECT 103.970 181.385 104.140 181.845 ;
        RECT 105.260 181.385 105.430 181.845 ;
        RECT 106.550 181.385 106.720 181.845 ;
        RECT 107.840 181.385 108.010 181.845 ;
        RECT 109.130 181.385 109.300 181.845 ;
        RECT 110.420 181.385 110.590 181.845 ;
        RECT 111.710 181.385 111.880 181.845 ;
        RECT 113.000 181.385 113.170 181.845 ;
        RECT 114.290 181.385 114.460 181.845 ;
        RECT 115.580 181.385 115.750 181.845 ;
        RECT 116.870 181.385 117.040 181.845 ;
        RECT 98.620 180.580 100.820 181.280 ;
        RECT 101.370 180.430 117.070 180.980 ;
        RECT 118.510 178.780 118.840 188.350 ;
        RECT 93.760 178.450 118.840 178.780 ;
        RECT 119.830 177.130 120.160 190.000 ;
        RECT 121.600 189.150 123.250 189.320 ;
        RECT 121.600 180.980 121.770 189.150 ;
        RECT 122.020 186.480 122.820 188.680 ;
        RECT 121.020 178.580 121.770 180.980 ;
        RECT 62.895 176.175 63.150 176.975 ;
        RECT 63.320 176.005 63.650 176.805 ;
        RECT 63.820 176.175 63.990 176.975 ;
        RECT 64.160 176.005 64.490 176.805 ;
        RECT 64.660 176.175 64.830 176.975 ;
        RECT 65.000 176.005 65.330 176.805 ;
        RECT 65.500 176.175 65.670 176.975 ;
        RECT 65.840 176.005 66.170 176.805 ;
        RECT 66.340 176.175 66.640 176.975 ;
        RECT 92.440 176.800 120.160 177.130 ;
        RECT 62.725 175.835 66.695 176.005 ;
        RECT 62.725 175.245 63.070 175.835 ;
        RECT 63.320 175.415 66.175 175.665 ;
        RECT 66.375 175.245 66.695 175.835 ;
        RECT 66.865 175.810 67.615 176.795 ;
        RECT 111.520 175.510 117.320 175.980 ;
        RECT 62.725 175.055 66.695 175.245 ;
        RECT 111.400 175.480 120.860 175.510 ;
        RECT 121.600 175.480 121.770 178.580 ;
        RECT 111.400 175.340 121.770 175.480 ;
        RECT 62.895 174.425 63.150 174.885 ;
        RECT 63.320 174.595 63.650 175.055 ;
        RECT 63.820 174.425 63.990 174.885 ;
        RECT 64.160 174.595 64.490 175.055 ;
        RECT 64.660 174.425 64.830 174.885 ;
        RECT 65.000 174.595 65.330 175.055 ;
        RECT 65.500 174.425 65.670 174.885 ;
        RECT 65.840 174.595 66.170 175.055 ;
        RECT 66.340 174.425 66.645 174.885 ;
        RECT 66.865 174.605 67.615 175.150 ;
        RECT 62.640 174.255 67.700 174.425 ;
        RECT 111.400 174.030 111.570 175.340 ;
        RECT 112.050 174.510 114.210 174.860 ;
        RECT 118.050 174.510 120.210 174.860 ;
        RECT 120.690 174.030 121.770 175.340 ;
        RECT 122.250 174.510 122.600 176.670 ;
        RECT 123.080 174.030 123.250 189.150 ;
        RECT 127.570 187.980 127.920 189.880 ;
        RECT 128.220 188.880 128.570 189.880 ;
        RECT 128.305 188.645 128.475 188.880 ;
        RECT 129.420 188.680 129.920 190.080 ;
        RECT 130.820 188.880 131.120 189.880 ;
        RECT 129.595 188.645 129.765 188.680 ;
        RECT 130.885 188.645 131.055 188.880 ;
        RECT 131.420 188.580 132.820 189.880 ;
        RECT 128.535 188.305 129.535 188.475 ;
        RECT 129.825 188.305 130.825 188.475 ;
        RECT 131.420 187.980 131.820 188.580 ;
        RECT 127.570 187.630 131.820 187.980 ;
        RECT 127.570 185.580 131.820 185.830 ;
        RECT 127.570 183.580 127.920 185.580 ;
        RECT 128.535 185.080 129.535 185.250 ;
        RECT 129.825 185.080 130.825 185.250 ;
        RECT 131.420 184.980 131.820 185.580 ;
        RECT 128.305 184.830 128.475 184.865 ;
        RECT 128.220 183.980 128.570 184.830 ;
        RECT 128.220 183.580 129.220 183.980 ;
        RECT 129.595 183.825 129.765 184.865 ;
        RECT 130.885 184.830 131.055 184.865 ;
        RECT 130.820 183.980 131.120 184.830 ;
        RECT 128.920 183.180 129.220 183.580 ;
        RECT 130.120 183.580 131.120 183.980 ;
        RECT 131.420 183.680 132.820 184.980 ;
        RECT 130.120 183.180 130.420 183.580 ;
        RECT 128.920 182.780 130.420 183.180 ;
        RECT 127.570 180.680 127.920 182.580 ;
        RECT 128.220 181.580 128.570 182.580 ;
        RECT 128.305 181.345 128.475 181.580 ;
        RECT 129.420 181.380 129.920 182.780 ;
        RECT 130.820 181.580 131.120 182.580 ;
        RECT 129.595 181.345 129.765 181.380 ;
        RECT 130.885 181.345 131.055 181.580 ;
        RECT 131.420 181.280 132.820 182.580 ;
        RECT 128.535 181.005 129.535 181.175 ;
        RECT 129.825 181.005 130.825 181.175 ;
        RECT 131.420 180.680 131.820 181.280 ;
        RECT 127.570 180.330 131.820 180.680 ;
        RECT 126.710 177.755 131.770 177.925 ;
        RECT 126.965 176.955 127.220 177.755 ;
        RECT 127.390 176.785 127.720 177.585 ;
        RECT 127.890 176.955 128.060 177.755 ;
        RECT 128.230 176.785 128.560 177.585 ;
        RECT 128.730 176.955 128.900 177.755 ;
        RECT 129.070 176.785 129.400 177.585 ;
        RECT 129.570 176.955 129.740 177.755 ;
        RECT 129.910 176.785 130.240 177.585 ;
        RECT 130.410 176.955 130.710 177.755 ;
        RECT 126.795 176.615 130.765 176.785 ;
        RECT 126.795 176.025 127.140 176.615 ;
        RECT 127.390 176.195 130.245 176.445 ;
        RECT 130.445 176.025 130.765 176.615 ;
        RECT 130.935 176.590 131.685 177.575 ;
        RECT 126.795 175.835 130.765 176.025 ;
        RECT 126.965 175.205 127.220 175.665 ;
        RECT 127.390 175.375 127.720 175.835 ;
        RECT 127.890 175.205 128.060 175.665 ;
        RECT 128.230 175.375 128.560 175.835 ;
        RECT 128.730 175.205 128.900 175.665 ;
        RECT 129.070 175.375 129.400 175.835 ;
        RECT 129.570 175.205 129.740 175.665 ;
        RECT 129.910 175.375 130.240 175.835 ;
        RECT 130.410 175.205 130.715 175.665 ;
        RECT 130.935 175.385 131.685 175.930 ;
        RECT 126.710 175.035 131.770 175.205 ;
        RECT 111.400 173.880 123.250 174.030 ;
        RECT 111.400 173.860 120.860 173.880 ;
        RECT 121.600 173.860 123.250 173.880 ;
        RECT 47.330 173.100 59.180 173.250 ;
        RECT 47.330 173.080 56.790 173.100 ;
        RECT 57.530 173.080 59.180 173.100 ;
        RECT 63.730 162.660 67.980 162.910 ;
        RECT 63.730 160.660 64.080 162.660 ;
        RECT 64.695 162.160 65.695 162.330 ;
        RECT 65.985 162.160 66.985 162.330 ;
        RECT 67.580 162.060 67.980 162.660 ;
        RECT 127.390 162.280 131.640 162.530 ;
        RECT 64.465 161.910 64.635 161.945 ;
        RECT 64.380 161.060 64.730 161.910 ;
        RECT 64.380 160.660 65.380 161.060 ;
        RECT 65.755 160.905 65.925 161.945 ;
        RECT 67.045 161.910 67.215 161.945 ;
        RECT 66.980 161.060 67.280 161.910 ;
        RECT 65.080 160.260 65.380 160.660 ;
        RECT 66.280 160.660 67.280 161.060 ;
        RECT 67.580 160.760 68.980 162.060 ;
        RECT 66.280 160.260 66.580 160.660 ;
        RECT 127.390 160.280 127.740 162.280 ;
        RECT 128.355 161.780 129.355 161.950 ;
        RECT 129.645 161.780 130.645 161.950 ;
        RECT 131.240 161.680 131.640 162.280 ;
        RECT 128.125 161.530 128.295 161.565 ;
        RECT 128.040 160.680 128.390 161.530 ;
        RECT 128.040 160.280 129.040 160.680 ;
        RECT 129.415 160.525 129.585 161.565 ;
        RECT 130.705 161.530 130.875 161.565 ;
        RECT 130.640 160.680 130.940 161.530 ;
        RECT 28.600 159.780 56.320 160.110 ;
        RECT 65.080 159.860 66.580 160.260 ;
        RECT 128.740 159.880 129.040 160.280 ;
        RECT 129.940 160.280 130.940 160.680 ;
        RECT 131.240 160.380 132.640 161.680 ;
        RECT 129.940 159.880 130.240 160.280 ;
        RECT 28.600 146.910 28.930 159.780 ;
        RECT 29.920 158.130 55.000 158.460 ;
        RECT 29.920 148.560 30.250 158.130 ;
        RECT 34.780 156.160 53.230 156.760 ;
        RECT 37.550 154.900 37.720 155.940 ;
        RECT 38.840 154.900 39.010 155.940 ;
        RECT 40.130 154.900 40.300 155.940 ;
        RECT 41.420 154.900 41.590 155.940 ;
        RECT 42.710 154.900 42.880 155.940 ;
        RECT 44.000 154.900 44.170 155.940 ;
        RECT 45.290 154.900 45.460 155.940 ;
        RECT 46.580 154.900 46.750 155.940 ;
        RECT 47.870 154.900 48.040 155.940 ;
        RECT 49.160 154.900 49.330 155.940 ;
        RECT 50.450 154.900 50.620 155.940 ;
        RECT 51.740 154.900 51.910 155.940 ;
        RECT 53.030 154.900 53.200 155.940 ;
        RECT 37.780 154.515 38.780 154.685 ;
        RECT 39.070 154.515 40.070 154.685 ;
        RECT 40.360 154.515 41.360 154.685 ;
        RECT 41.650 154.515 42.650 154.685 ;
        RECT 42.940 154.515 43.940 154.685 ;
        RECT 44.230 154.515 45.230 154.685 ;
        RECT 45.520 154.515 46.520 154.685 ;
        RECT 46.810 154.515 47.810 154.685 ;
        RECT 48.100 154.515 49.100 154.685 ;
        RECT 49.390 154.515 50.390 154.685 ;
        RECT 50.680 154.515 51.680 154.685 ;
        RECT 51.970 154.515 52.970 154.685 ;
        RECT 39.070 153.975 40.070 154.145 ;
        RECT 42.940 153.975 43.940 154.145 ;
        RECT 44.230 153.975 45.230 154.145 ;
        RECT 48.100 153.975 49.100 154.145 ;
        RECT 49.390 153.975 50.390 154.145 ;
        RECT 37.550 152.765 37.720 153.805 ;
        RECT 38.840 152.765 39.010 153.805 ;
        RECT 40.130 152.765 40.300 153.805 ;
        RECT 41.420 152.765 41.590 153.805 ;
        RECT 42.710 152.765 42.880 153.805 ;
        RECT 44.000 152.765 44.170 153.805 ;
        RECT 45.290 152.765 45.460 153.805 ;
        RECT 46.580 152.765 46.750 153.805 ;
        RECT 47.870 152.765 48.040 153.805 ;
        RECT 49.160 152.765 49.330 153.805 ;
        RECT 50.450 152.765 50.620 153.805 ;
        RECT 51.740 152.765 51.910 153.805 ;
        RECT 53.030 152.765 53.200 153.805 ;
        RECT 37.780 152.425 38.780 152.595 ;
        RECT 40.360 152.425 41.360 152.595 ;
        RECT 41.650 152.425 42.650 152.595 ;
        RECT 45.520 152.425 46.520 152.595 ;
        RECT 46.810 152.425 47.810 152.595 ;
        RECT 50.680 152.425 51.680 152.595 ;
        RECT 51.970 152.425 52.970 152.595 ;
        RECT 37.780 151.795 38.780 151.965 ;
        RECT 39.070 151.795 40.070 151.965 ;
        RECT 40.360 151.795 41.360 151.965 ;
        RECT 41.650 151.795 42.650 151.965 ;
        RECT 42.940 151.795 43.940 151.965 ;
        RECT 44.230 151.795 45.230 151.965 ;
        RECT 45.520 151.795 46.520 151.965 ;
        RECT 46.810 151.795 47.810 151.965 ;
        RECT 48.100 151.795 49.100 151.965 ;
        RECT 49.390 151.795 50.390 151.965 ;
        RECT 50.680 151.795 51.680 151.965 ;
        RECT 51.970 151.795 52.970 151.965 ;
        RECT 37.550 151.165 37.720 151.625 ;
        RECT 38.840 151.165 39.010 151.625 ;
        RECT 40.130 151.165 40.300 151.625 ;
        RECT 41.420 151.165 41.590 151.625 ;
        RECT 42.710 151.165 42.880 151.625 ;
        RECT 44.000 151.165 44.170 151.625 ;
        RECT 45.290 151.165 45.460 151.625 ;
        RECT 46.580 151.165 46.750 151.625 ;
        RECT 47.870 151.165 48.040 151.625 ;
        RECT 49.160 151.165 49.330 151.625 ;
        RECT 50.450 151.165 50.620 151.625 ;
        RECT 51.740 151.165 51.910 151.625 ;
        RECT 53.030 151.165 53.200 151.625 ;
        RECT 34.780 150.360 36.980 151.060 ;
        RECT 37.530 150.210 53.230 150.760 ;
        RECT 54.670 148.560 55.000 158.130 ;
        RECT 29.920 148.230 55.000 148.560 ;
        RECT 55.990 146.910 56.320 159.780 ;
        RECT 57.760 158.930 59.410 159.100 ;
        RECT 57.760 150.760 57.930 158.930 ;
        RECT 58.180 156.260 58.980 158.460 ;
        RECT 57.180 148.360 57.930 150.760 ;
        RECT 28.600 146.580 56.320 146.910 ;
        RECT 47.680 145.290 53.480 145.760 ;
        RECT 47.560 145.260 57.020 145.290 ;
        RECT 57.760 145.260 57.930 148.360 ;
        RECT 47.560 145.120 57.930 145.260 ;
        RECT 47.560 143.810 47.730 145.120 ;
        RECT 48.210 144.290 50.370 144.640 ;
        RECT 54.210 144.290 56.370 144.640 ;
        RECT 56.850 143.810 57.930 145.120 ;
        RECT 58.410 144.290 58.760 146.450 ;
        RECT 59.240 143.810 59.410 158.930 ;
        RECT 63.730 157.760 64.080 159.660 ;
        RECT 64.380 158.660 64.730 159.660 ;
        RECT 64.465 158.425 64.635 158.660 ;
        RECT 65.580 158.460 66.080 159.860 ;
        RECT 66.980 158.660 67.280 159.660 ;
        RECT 65.755 158.425 65.925 158.460 ;
        RECT 67.045 158.425 67.215 158.660 ;
        RECT 67.580 158.360 68.980 159.660 ;
        RECT 92.260 159.400 119.980 159.730 ;
        RECT 128.740 159.480 130.240 159.880 ;
        RECT 64.695 158.085 65.695 158.255 ;
        RECT 65.985 158.085 66.985 158.255 ;
        RECT 67.580 157.760 67.980 158.360 ;
        RECT 63.730 157.410 67.980 157.760 ;
        RECT 63.730 155.360 67.980 155.610 ;
        RECT 63.730 153.360 64.080 155.360 ;
        RECT 64.695 154.860 65.695 155.030 ;
        RECT 65.985 154.860 66.985 155.030 ;
        RECT 67.580 154.760 67.980 155.360 ;
        RECT 64.465 154.610 64.635 154.645 ;
        RECT 64.380 153.760 64.730 154.610 ;
        RECT 64.380 153.360 65.380 153.760 ;
        RECT 65.755 153.605 65.925 154.645 ;
        RECT 67.045 154.610 67.215 154.645 ;
        RECT 66.980 153.760 67.280 154.610 ;
        RECT 65.080 152.960 65.380 153.360 ;
        RECT 66.280 153.360 67.280 153.760 ;
        RECT 67.580 153.460 68.980 154.760 ;
        RECT 66.280 152.960 66.580 153.360 ;
        RECT 65.080 152.560 66.580 152.960 ;
        RECT 63.730 150.460 64.080 152.360 ;
        RECT 64.380 151.360 64.730 152.360 ;
        RECT 64.465 151.125 64.635 151.360 ;
        RECT 65.580 151.160 66.080 152.560 ;
        RECT 66.980 151.360 67.280 152.360 ;
        RECT 65.755 151.125 65.925 151.160 ;
        RECT 67.045 151.125 67.215 151.360 ;
        RECT 67.580 151.060 68.980 152.360 ;
        RECT 64.695 150.785 65.695 150.955 ;
        RECT 65.985 150.785 66.985 150.955 ;
        RECT 67.580 150.460 67.980 151.060 ;
        RECT 63.730 150.110 67.980 150.460 ;
        RECT 62.870 147.535 67.930 147.705 ;
        RECT 63.125 146.735 63.380 147.535 ;
        RECT 63.550 146.565 63.880 147.365 ;
        RECT 64.050 146.735 64.220 147.535 ;
        RECT 64.390 146.565 64.720 147.365 ;
        RECT 64.890 146.735 65.060 147.535 ;
        RECT 65.230 146.565 65.560 147.365 ;
        RECT 65.730 146.735 65.900 147.535 ;
        RECT 66.070 146.565 66.400 147.365 ;
        RECT 66.570 146.735 66.870 147.535 ;
        RECT 62.955 146.395 66.925 146.565 ;
        RECT 62.955 145.805 63.300 146.395 ;
        RECT 63.550 145.975 66.405 146.225 ;
        RECT 66.605 145.805 66.925 146.395 ;
        RECT 67.095 146.370 67.845 147.355 ;
        RECT 92.260 146.530 92.590 159.400 ;
        RECT 93.580 157.750 118.660 158.080 ;
        RECT 93.580 148.180 93.910 157.750 ;
        RECT 98.440 155.780 116.890 156.380 ;
        RECT 101.210 154.520 101.380 155.560 ;
        RECT 102.500 154.520 102.670 155.560 ;
        RECT 103.790 154.520 103.960 155.560 ;
        RECT 105.080 154.520 105.250 155.560 ;
        RECT 106.370 154.520 106.540 155.560 ;
        RECT 107.660 154.520 107.830 155.560 ;
        RECT 108.950 154.520 109.120 155.560 ;
        RECT 110.240 154.520 110.410 155.560 ;
        RECT 111.530 154.520 111.700 155.560 ;
        RECT 112.820 154.520 112.990 155.560 ;
        RECT 114.110 154.520 114.280 155.560 ;
        RECT 115.400 154.520 115.570 155.560 ;
        RECT 116.690 154.520 116.860 155.560 ;
        RECT 101.440 154.135 102.440 154.305 ;
        RECT 102.730 154.135 103.730 154.305 ;
        RECT 104.020 154.135 105.020 154.305 ;
        RECT 105.310 154.135 106.310 154.305 ;
        RECT 106.600 154.135 107.600 154.305 ;
        RECT 107.890 154.135 108.890 154.305 ;
        RECT 109.180 154.135 110.180 154.305 ;
        RECT 110.470 154.135 111.470 154.305 ;
        RECT 111.760 154.135 112.760 154.305 ;
        RECT 113.050 154.135 114.050 154.305 ;
        RECT 114.340 154.135 115.340 154.305 ;
        RECT 115.630 154.135 116.630 154.305 ;
        RECT 102.730 153.595 103.730 153.765 ;
        RECT 106.600 153.595 107.600 153.765 ;
        RECT 107.890 153.595 108.890 153.765 ;
        RECT 111.760 153.595 112.760 153.765 ;
        RECT 113.050 153.595 114.050 153.765 ;
        RECT 101.210 152.385 101.380 153.425 ;
        RECT 102.500 152.385 102.670 153.425 ;
        RECT 103.790 152.385 103.960 153.425 ;
        RECT 105.080 152.385 105.250 153.425 ;
        RECT 106.370 152.385 106.540 153.425 ;
        RECT 107.660 152.385 107.830 153.425 ;
        RECT 108.950 152.385 109.120 153.425 ;
        RECT 110.240 152.385 110.410 153.425 ;
        RECT 111.530 152.385 111.700 153.425 ;
        RECT 112.820 152.385 112.990 153.425 ;
        RECT 114.110 152.385 114.280 153.425 ;
        RECT 115.400 152.385 115.570 153.425 ;
        RECT 116.690 152.385 116.860 153.425 ;
        RECT 101.440 152.045 102.440 152.215 ;
        RECT 104.020 152.045 105.020 152.215 ;
        RECT 105.310 152.045 106.310 152.215 ;
        RECT 109.180 152.045 110.180 152.215 ;
        RECT 110.470 152.045 111.470 152.215 ;
        RECT 114.340 152.045 115.340 152.215 ;
        RECT 115.630 152.045 116.630 152.215 ;
        RECT 101.440 151.415 102.440 151.585 ;
        RECT 102.730 151.415 103.730 151.585 ;
        RECT 104.020 151.415 105.020 151.585 ;
        RECT 105.310 151.415 106.310 151.585 ;
        RECT 106.600 151.415 107.600 151.585 ;
        RECT 107.890 151.415 108.890 151.585 ;
        RECT 109.180 151.415 110.180 151.585 ;
        RECT 110.470 151.415 111.470 151.585 ;
        RECT 111.760 151.415 112.760 151.585 ;
        RECT 113.050 151.415 114.050 151.585 ;
        RECT 114.340 151.415 115.340 151.585 ;
        RECT 115.630 151.415 116.630 151.585 ;
        RECT 101.210 150.785 101.380 151.245 ;
        RECT 102.500 150.785 102.670 151.245 ;
        RECT 103.790 150.785 103.960 151.245 ;
        RECT 105.080 150.785 105.250 151.245 ;
        RECT 106.370 150.785 106.540 151.245 ;
        RECT 107.660 150.785 107.830 151.245 ;
        RECT 108.950 150.785 109.120 151.245 ;
        RECT 110.240 150.785 110.410 151.245 ;
        RECT 111.530 150.785 111.700 151.245 ;
        RECT 112.820 150.785 112.990 151.245 ;
        RECT 114.110 150.785 114.280 151.245 ;
        RECT 115.400 150.785 115.570 151.245 ;
        RECT 116.690 150.785 116.860 151.245 ;
        RECT 98.440 149.980 100.640 150.680 ;
        RECT 101.190 149.830 116.890 150.380 ;
        RECT 118.330 148.180 118.660 157.750 ;
        RECT 93.580 147.850 118.660 148.180 ;
        RECT 119.650 146.530 119.980 159.400 ;
        RECT 121.420 158.550 123.070 158.720 ;
        RECT 121.420 150.380 121.590 158.550 ;
        RECT 121.840 155.880 122.640 158.080 ;
        RECT 120.840 147.980 121.590 150.380 ;
        RECT 92.260 146.200 119.980 146.530 ;
        RECT 62.955 145.615 66.925 145.805 ;
        RECT 63.125 144.985 63.380 145.445 ;
        RECT 63.550 145.155 63.880 145.615 ;
        RECT 64.050 144.985 64.220 145.445 ;
        RECT 64.390 145.155 64.720 145.615 ;
        RECT 64.890 144.985 65.060 145.445 ;
        RECT 65.230 145.155 65.560 145.615 ;
        RECT 65.730 144.985 65.900 145.445 ;
        RECT 66.070 145.155 66.400 145.615 ;
        RECT 66.570 144.985 66.875 145.445 ;
        RECT 67.095 145.165 67.845 145.710 ;
        RECT 62.870 144.815 67.930 144.985 ;
        RECT 111.340 144.910 117.140 145.380 ;
        RECT 111.220 144.880 120.680 144.910 ;
        RECT 121.420 144.880 121.590 147.980 ;
        RECT 47.560 143.660 59.410 143.810 ;
        RECT 47.560 143.640 57.020 143.660 ;
        RECT 57.760 143.640 59.410 143.660 ;
        RECT 111.220 144.740 121.590 144.880 ;
        RECT 111.220 143.430 111.390 144.740 ;
        RECT 111.870 143.910 114.030 144.260 ;
        RECT 117.870 143.910 120.030 144.260 ;
        RECT 120.510 143.430 121.590 144.740 ;
        RECT 122.070 143.910 122.420 146.070 ;
        RECT 122.900 143.430 123.070 158.550 ;
        RECT 127.390 157.380 127.740 159.280 ;
        RECT 128.040 158.280 128.390 159.280 ;
        RECT 128.125 158.045 128.295 158.280 ;
        RECT 129.240 158.080 129.740 159.480 ;
        RECT 130.640 158.280 130.940 159.280 ;
        RECT 129.415 158.045 129.585 158.080 ;
        RECT 130.705 158.045 130.875 158.280 ;
        RECT 131.240 157.980 132.640 159.280 ;
        RECT 128.355 157.705 129.355 157.875 ;
        RECT 129.645 157.705 130.645 157.875 ;
        RECT 131.240 157.380 131.640 157.980 ;
        RECT 127.390 157.030 131.640 157.380 ;
        RECT 127.390 154.980 131.640 155.230 ;
        RECT 127.390 152.980 127.740 154.980 ;
        RECT 128.355 154.480 129.355 154.650 ;
        RECT 129.645 154.480 130.645 154.650 ;
        RECT 131.240 154.380 131.640 154.980 ;
        RECT 128.125 154.230 128.295 154.265 ;
        RECT 128.040 153.380 128.390 154.230 ;
        RECT 128.040 152.980 129.040 153.380 ;
        RECT 129.415 153.225 129.585 154.265 ;
        RECT 130.705 154.230 130.875 154.265 ;
        RECT 130.640 153.380 130.940 154.230 ;
        RECT 128.740 152.580 129.040 152.980 ;
        RECT 129.940 152.980 130.940 153.380 ;
        RECT 131.240 153.080 132.640 154.380 ;
        RECT 129.940 152.580 130.240 152.980 ;
        RECT 128.740 152.180 130.240 152.580 ;
        RECT 127.390 150.080 127.740 151.980 ;
        RECT 128.040 150.980 128.390 151.980 ;
        RECT 128.125 150.745 128.295 150.980 ;
        RECT 129.240 150.780 129.740 152.180 ;
        RECT 130.640 150.980 130.940 151.980 ;
        RECT 129.415 150.745 129.585 150.780 ;
        RECT 130.705 150.745 130.875 150.980 ;
        RECT 131.240 150.680 132.640 151.980 ;
        RECT 128.355 150.405 129.355 150.575 ;
        RECT 129.645 150.405 130.645 150.575 ;
        RECT 131.240 150.080 131.640 150.680 ;
        RECT 127.390 149.730 131.640 150.080 ;
        RECT 126.530 147.155 131.590 147.325 ;
        RECT 126.785 146.355 127.040 147.155 ;
        RECT 127.210 146.185 127.540 146.985 ;
        RECT 127.710 146.355 127.880 147.155 ;
        RECT 128.050 146.185 128.380 146.985 ;
        RECT 128.550 146.355 128.720 147.155 ;
        RECT 128.890 146.185 129.220 146.985 ;
        RECT 129.390 146.355 129.560 147.155 ;
        RECT 129.730 146.185 130.060 146.985 ;
        RECT 130.230 146.355 130.530 147.155 ;
        RECT 126.615 146.015 130.585 146.185 ;
        RECT 126.615 145.425 126.960 146.015 ;
        RECT 127.210 145.595 130.065 145.845 ;
        RECT 130.265 145.425 130.585 146.015 ;
        RECT 130.755 145.990 131.505 146.975 ;
        RECT 126.615 145.235 130.585 145.425 ;
        RECT 126.785 144.605 127.040 145.065 ;
        RECT 127.210 144.775 127.540 145.235 ;
        RECT 127.710 144.605 127.880 145.065 ;
        RECT 128.050 144.775 128.380 145.235 ;
        RECT 128.550 144.605 128.720 145.065 ;
        RECT 128.890 144.775 129.220 145.235 ;
        RECT 129.390 144.605 129.560 145.065 ;
        RECT 129.730 144.775 130.060 145.235 ;
        RECT 130.230 144.605 130.535 145.065 ;
        RECT 130.755 144.785 131.505 145.330 ;
        RECT 126.530 144.435 131.590 144.605 ;
        RECT 111.220 143.280 123.070 143.430 ;
        RECT 111.220 143.260 120.680 143.280 ;
        RECT 121.420 143.260 123.070 143.280 ;
        RECT 64.330 129.140 68.580 129.390 ;
        RECT 64.330 127.140 64.680 129.140 ;
        RECT 65.295 128.640 66.295 128.810 ;
        RECT 66.585 128.640 67.585 128.810 ;
        RECT 68.180 128.540 68.580 129.140 ;
        RECT 65.065 128.390 65.235 128.425 ;
        RECT 64.980 127.540 65.330 128.390 ;
        RECT 64.980 127.140 65.980 127.540 ;
        RECT 66.355 127.385 66.525 128.425 ;
        RECT 67.645 128.390 67.815 128.425 ;
        RECT 67.580 127.540 67.880 128.390 ;
        RECT 65.680 126.740 65.980 127.140 ;
        RECT 66.880 127.140 67.880 127.540 ;
        RECT 68.180 127.240 69.580 128.540 ;
        RECT 127.870 128.490 132.120 128.740 ;
        RECT 66.880 126.740 67.180 127.140 ;
        RECT 29.200 126.260 56.920 126.590 ;
        RECT 65.680 126.340 67.180 126.740 ;
        RECT 127.870 126.490 128.220 128.490 ;
        RECT 128.835 127.990 129.835 128.160 ;
        RECT 130.125 127.990 131.125 128.160 ;
        RECT 131.720 127.890 132.120 128.490 ;
        RECT 128.605 127.740 128.775 127.775 ;
        RECT 128.520 126.890 128.870 127.740 ;
        RECT 128.520 126.490 129.520 126.890 ;
        RECT 129.895 126.735 130.065 127.775 ;
        RECT 131.185 127.740 131.355 127.775 ;
        RECT 131.120 126.890 131.420 127.740 ;
        RECT 29.200 113.390 29.530 126.260 ;
        RECT 30.520 124.610 55.600 124.940 ;
        RECT 30.520 115.040 30.850 124.610 ;
        RECT 35.380 122.640 53.830 123.240 ;
        RECT 38.150 121.380 38.320 122.420 ;
        RECT 39.440 121.380 39.610 122.420 ;
        RECT 40.730 121.380 40.900 122.420 ;
        RECT 42.020 121.380 42.190 122.420 ;
        RECT 43.310 121.380 43.480 122.420 ;
        RECT 44.600 121.380 44.770 122.420 ;
        RECT 45.890 121.380 46.060 122.420 ;
        RECT 47.180 121.380 47.350 122.420 ;
        RECT 48.470 121.380 48.640 122.420 ;
        RECT 49.760 121.380 49.930 122.420 ;
        RECT 51.050 121.380 51.220 122.420 ;
        RECT 52.340 121.380 52.510 122.420 ;
        RECT 53.630 121.380 53.800 122.420 ;
        RECT 38.380 120.995 39.380 121.165 ;
        RECT 39.670 120.995 40.670 121.165 ;
        RECT 40.960 120.995 41.960 121.165 ;
        RECT 42.250 120.995 43.250 121.165 ;
        RECT 43.540 120.995 44.540 121.165 ;
        RECT 44.830 120.995 45.830 121.165 ;
        RECT 46.120 120.995 47.120 121.165 ;
        RECT 47.410 120.995 48.410 121.165 ;
        RECT 48.700 120.995 49.700 121.165 ;
        RECT 49.990 120.995 50.990 121.165 ;
        RECT 51.280 120.995 52.280 121.165 ;
        RECT 52.570 120.995 53.570 121.165 ;
        RECT 39.670 120.455 40.670 120.625 ;
        RECT 43.540 120.455 44.540 120.625 ;
        RECT 44.830 120.455 45.830 120.625 ;
        RECT 48.700 120.455 49.700 120.625 ;
        RECT 49.990 120.455 50.990 120.625 ;
        RECT 38.150 119.245 38.320 120.285 ;
        RECT 39.440 119.245 39.610 120.285 ;
        RECT 40.730 119.245 40.900 120.285 ;
        RECT 42.020 119.245 42.190 120.285 ;
        RECT 43.310 119.245 43.480 120.285 ;
        RECT 44.600 119.245 44.770 120.285 ;
        RECT 45.890 119.245 46.060 120.285 ;
        RECT 47.180 119.245 47.350 120.285 ;
        RECT 48.470 119.245 48.640 120.285 ;
        RECT 49.760 119.245 49.930 120.285 ;
        RECT 51.050 119.245 51.220 120.285 ;
        RECT 52.340 119.245 52.510 120.285 ;
        RECT 53.630 119.245 53.800 120.285 ;
        RECT 38.380 118.905 39.380 119.075 ;
        RECT 40.960 118.905 41.960 119.075 ;
        RECT 42.250 118.905 43.250 119.075 ;
        RECT 46.120 118.905 47.120 119.075 ;
        RECT 47.410 118.905 48.410 119.075 ;
        RECT 51.280 118.905 52.280 119.075 ;
        RECT 52.570 118.905 53.570 119.075 ;
        RECT 38.380 118.275 39.380 118.445 ;
        RECT 39.670 118.275 40.670 118.445 ;
        RECT 40.960 118.275 41.960 118.445 ;
        RECT 42.250 118.275 43.250 118.445 ;
        RECT 43.540 118.275 44.540 118.445 ;
        RECT 44.830 118.275 45.830 118.445 ;
        RECT 46.120 118.275 47.120 118.445 ;
        RECT 47.410 118.275 48.410 118.445 ;
        RECT 48.700 118.275 49.700 118.445 ;
        RECT 49.990 118.275 50.990 118.445 ;
        RECT 51.280 118.275 52.280 118.445 ;
        RECT 52.570 118.275 53.570 118.445 ;
        RECT 38.150 117.645 38.320 118.105 ;
        RECT 39.440 117.645 39.610 118.105 ;
        RECT 40.730 117.645 40.900 118.105 ;
        RECT 42.020 117.645 42.190 118.105 ;
        RECT 43.310 117.645 43.480 118.105 ;
        RECT 44.600 117.645 44.770 118.105 ;
        RECT 45.890 117.645 46.060 118.105 ;
        RECT 47.180 117.645 47.350 118.105 ;
        RECT 48.470 117.645 48.640 118.105 ;
        RECT 49.760 117.645 49.930 118.105 ;
        RECT 51.050 117.645 51.220 118.105 ;
        RECT 52.340 117.645 52.510 118.105 ;
        RECT 53.630 117.645 53.800 118.105 ;
        RECT 35.380 116.840 37.580 117.540 ;
        RECT 38.130 116.690 53.830 117.240 ;
        RECT 55.270 115.040 55.600 124.610 ;
        RECT 30.520 114.710 55.600 115.040 ;
        RECT 56.590 113.390 56.920 126.260 ;
        RECT 58.360 125.410 60.010 125.580 ;
        RECT 58.360 117.240 58.530 125.410 ;
        RECT 58.780 122.740 59.580 124.940 ;
        RECT 57.780 114.840 58.530 117.240 ;
        RECT 29.200 113.060 56.920 113.390 ;
        RECT 48.280 111.770 54.080 112.240 ;
        RECT 48.160 111.740 57.620 111.770 ;
        RECT 58.360 111.740 58.530 114.840 ;
        RECT 48.160 111.600 58.530 111.740 ;
        RECT 48.160 110.290 48.330 111.600 ;
        RECT 48.810 110.770 50.970 111.120 ;
        RECT 54.810 110.770 56.970 111.120 ;
        RECT 57.450 110.290 58.530 111.600 ;
        RECT 59.010 110.770 59.360 112.930 ;
        RECT 59.840 110.290 60.010 125.410 ;
        RECT 64.330 124.240 64.680 126.140 ;
        RECT 64.980 125.140 65.330 126.140 ;
        RECT 65.065 124.905 65.235 125.140 ;
        RECT 66.180 124.940 66.680 126.340 ;
        RECT 67.580 125.140 67.880 126.140 ;
        RECT 66.355 124.905 66.525 124.940 ;
        RECT 67.645 124.905 67.815 125.140 ;
        RECT 68.180 124.840 69.580 126.140 ;
        RECT 129.220 126.090 129.520 126.490 ;
        RECT 130.420 126.490 131.420 126.890 ;
        RECT 131.720 126.590 133.120 127.890 ;
        RECT 130.420 126.090 130.720 126.490 ;
        RECT 92.740 125.610 120.460 125.940 ;
        RECT 129.220 125.690 130.720 126.090 ;
        RECT 65.295 124.565 66.295 124.735 ;
        RECT 66.585 124.565 67.585 124.735 ;
        RECT 68.180 124.240 68.580 124.840 ;
        RECT 64.330 123.890 68.580 124.240 ;
        RECT 64.330 121.840 68.580 122.090 ;
        RECT 64.330 119.840 64.680 121.840 ;
        RECT 65.295 121.340 66.295 121.510 ;
        RECT 66.585 121.340 67.585 121.510 ;
        RECT 68.180 121.240 68.580 121.840 ;
        RECT 65.065 121.090 65.235 121.125 ;
        RECT 64.980 120.240 65.330 121.090 ;
        RECT 64.980 119.840 65.980 120.240 ;
        RECT 66.355 120.085 66.525 121.125 ;
        RECT 67.645 121.090 67.815 121.125 ;
        RECT 67.580 120.240 67.880 121.090 ;
        RECT 65.680 119.440 65.980 119.840 ;
        RECT 66.880 119.840 67.880 120.240 ;
        RECT 68.180 119.940 69.580 121.240 ;
        RECT 66.880 119.440 67.180 119.840 ;
        RECT 65.680 119.040 67.180 119.440 ;
        RECT 64.330 116.940 64.680 118.840 ;
        RECT 64.980 117.840 65.330 118.840 ;
        RECT 65.065 117.605 65.235 117.840 ;
        RECT 66.180 117.640 66.680 119.040 ;
        RECT 67.580 117.840 67.880 118.840 ;
        RECT 66.355 117.605 66.525 117.640 ;
        RECT 67.645 117.605 67.815 117.840 ;
        RECT 68.180 117.540 69.580 118.840 ;
        RECT 65.295 117.265 66.295 117.435 ;
        RECT 66.585 117.265 67.585 117.435 ;
        RECT 68.180 116.940 68.580 117.540 ;
        RECT 64.330 116.590 68.580 116.940 ;
        RECT 63.470 114.015 68.530 114.185 ;
        RECT 63.725 113.215 63.980 114.015 ;
        RECT 64.150 113.045 64.480 113.845 ;
        RECT 64.650 113.215 64.820 114.015 ;
        RECT 64.990 113.045 65.320 113.845 ;
        RECT 65.490 113.215 65.660 114.015 ;
        RECT 65.830 113.045 66.160 113.845 ;
        RECT 66.330 113.215 66.500 114.015 ;
        RECT 66.670 113.045 67.000 113.845 ;
        RECT 67.170 113.215 67.470 114.015 ;
        RECT 63.555 112.875 67.525 113.045 ;
        RECT 63.555 112.285 63.900 112.875 ;
        RECT 64.150 112.455 67.005 112.705 ;
        RECT 67.205 112.285 67.525 112.875 ;
        RECT 67.695 112.850 68.445 113.835 ;
        RECT 92.740 112.740 93.070 125.610 ;
        RECT 94.060 123.960 119.140 124.290 ;
        RECT 94.060 114.390 94.390 123.960 ;
        RECT 98.920 121.990 117.370 122.590 ;
        RECT 101.690 120.730 101.860 121.770 ;
        RECT 102.980 120.730 103.150 121.770 ;
        RECT 104.270 120.730 104.440 121.770 ;
        RECT 105.560 120.730 105.730 121.770 ;
        RECT 106.850 120.730 107.020 121.770 ;
        RECT 108.140 120.730 108.310 121.770 ;
        RECT 109.430 120.730 109.600 121.770 ;
        RECT 110.720 120.730 110.890 121.770 ;
        RECT 112.010 120.730 112.180 121.770 ;
        RECT 113.300 120.730 113.470 121.770 ;
        RECT 114.590 120.730 114.760 121.770 ;
        RECT 115.880 120.730 116.050 121.770 ;
        RECT 117.170 120.730 117.340 121.770 ;
        RECT 101.920 120.345 102.920 120.515 ;
        RECT 103.210 120.345 104.210 120.515 ;
        RECT 104.500 120.345 105.500 120.515 ;
        RECT 105.790 120.345 106.790 120.515 ;
        RECT 107.080 120.345 108.080 120.515 ;
        RECT 108.370 120.345 109.370 120.515 ;
        RECT 109.660 120.345 110.660 120.515 ;
        RECT 110.950 120.345 111.950 120.515 ;
        RECT 112.240 120.345 113.240 120.515 ;
        RECT 113.530 120.345 114.530 120.515 ;
        RECT 114.820 120.345 115.820 120.515 ;
        RECT 116.110 120.345 117.110 120.515 ;
        RECT 103.210 119.805 104.210 119.975 ;
        RECT 107.080 119.805 108.080 119.975 ;
        RECT 108.370 119.805 109.370 119.975 ;
        RECT 112.240 119.805 113.240 119.975 ;
        RECT 113.530 119.805 114.530 119.975 ;
        RECT 101.690 118.595 101.860 119.635 ;
        RECT 102.980 118.595 103.150 119.635 ;
        RECT 104.270 118.595 104.440 119.635 ;
        RECT 105.560 118.595 105.730 119.635 ;
        RECT 106.850 118.595 107.020 119.635 ;
        RECT 108.140 118.595 108.310 119.635 ;
        RECT 109.430 118.595 109.600 119.635 ;
        RECT 110.720 118.595 110.890 119.635 ;
        RECT 112.010 118.595 112.180 119.635 ;
        RECT 113.300 118.595 113.470 119.635 ;
        RECT 114.590 118.595 114.760 119.635 ;
        RECT 115.880 118.595 116.050 119.635 ;
        RECT 117.170 118.595 117.340 119.635 ;
        RECT 101.920 118.255 102.920 118.425 ;
        RECT 104.500 118.255 105.500 118.425 ;
        RECT 105.790 118.255 106.790 118.425 ;
        RECT 109.660 118.255 110.660 118.425 ;
        RECT 110.950 118.255 111.950 118.425 ;
        RECT 114.820 118.255 115.820 118.425 ;
        RECT 116.110 118.255 117.110 118.425 ;
        RECT 101.920 117.625 102.920 117.795 ;
        RECT 103.210 117.625 104.210 117.795 ;
        RECT 104.500 117.625 105.500 117.795 ;
        RECT 105.790 117.625 106.790 117.795 ;
        RECT 107.080 117.625 108.080 117.795 ;
        RECT 108.370 117.625 109.370 117.795 ;
        RECT 109.660 117.625 110.660 117.795 ;
        RECT 110.950 117.625 111.950 117.795 ;
        RECT 112.240 117.625 113.240 117.795 ;
        RECT 113.530 117.625 114.530 117.795 ;
        RECT 114.820 117.625 115.820 117.795 ;
        RECT 116.110 117.625 117.110 117.795 ;
        RECT 101.690 116.995 101.860 117.455 ;
        RECT 102.980 116.995 103.150 117.455 ;
        RECT 104.270 116.995 104.440 117.455 ;
        RECT 105.560 116.995 105.730 117.455 ;
        RECT 106.850 116.995 107.020 117.455 ;
        RECT 108.140 116.995 108.310 117.455 ;
        RECT 109.430 116.995 109.600 117.455 ;
        RECT 110.720 116.995 110.890 117.455 ;
        RECT 112.010 116.995 112.180 117.455 ;
        RECT 113.300 116.995 113.470 117.455 ;
        RECT 114.590 116.995 114.760 117.455 ;
        RECT 115.880 116.995 116.050 117.455 ;
        RECT 117.170 116.995 117.340 117.455 ;
        RECT 98.920 116.190 101.120 116.890 ;
        RECT 101.670 116.040 117.370 116.590 ;
        RECT 118.810 114.390 119.140 123.960 ;
        RECT 94.060 114.060 119.140 114.390 ;
        RECT 120.130 112.740 120.460 125.610 ;
        RECT 121.900 124.760 123.550 124.930 ;
        RECT 121.900 116.590 122.070 124.760 ;
        RECT 122.320 122.090 123.120 124.290 ;
        RECT 121.320 114.190 122.070 116.590 ;
        RECT 92.740 112.410 120.460 112.740 ;
        RECT 63.555 112.095 67.525 112.285 ;
        RECT 63.725 111.465 63.980 111.925 ;
        RECT 64.150 111.635 64.480 112.095 ;
        RECT 64.650 111.465 64.820 111.925 ;
        RECT 64.990 111.635 65.320 112.095 ;
        RECT 65.490 111.465 65.660 111.925 ;
        RECT 65.830 111.635 66.160 112.095 ;
        RECT 66.330 111.465 66.500 111.925 ;
        RECT 66.670 111.635 67.000 112.095 ;
        RECT 67.170 111.465 67.475 111.925 ;
        RECT 67.695 111.645 68.445 112.190 ;
        RECT 63.470 111.295 68.530 111.465 ;
        RECT 111.820 111.120 117.620 111.590 ;
        RECT 48.160 110.140 60.010 110.290 ;
        RECT 48.160 110.120 57.620 110.140 ;
        RECT 58.360 110.120 60.010 110.140 ;
        RECT 111.700 111.090 121.160 111.120 ;
        RECT 121.900 111.090 122.070 114.190 ;
        RECT 111.700 110.950 122.070 111.090 ;
        RECT 111.700 109.640 111.870 110.950 ;
        RECT 112.350 110.120 114.510 110.470 ;
        RECT 118.350 110.120 120.510 110.470 ;
        RECT 120.990 109.640 122.070 110.950 ;
        RECT 122.550 110.120 122.900 112.280 ;
        RECT 123.380 109.640 123.550 124.760 ;
        RECT 127.870 123.590 128.220 125.490 ;
        RECT 128.520 124.490 128.870 125.490 ;
        RECT 128.605 124.255 128.775 124.490 ;
        RECT 129.720 124.290 130.220 125.690 ;
        RECT 131.120 124.490 131.420 125.490 ;
        RECT 129.895 124.255 130.065 124.290 ;
        RECT 131.185 124.255 131.355 124.490 ;
        RECT 131.720 124.190 133.120 125.490 ;
        RECT 128.835 123.915 129.835 124.085 ;
        RECT 130.125 123.915 131.125 124.085 ;
        RECT 131.720 123.590 132.120 124.190 ;
        RECT 127.870 123.240 132.120 123.590 ;
        RECT 127.870 121.190 132.120 121.440 ;
        RECT 127.870 119.190 128.220 121.190 ;
        RECT 128.835 120.690 129.835 120.860 ;
        RECT 130.125 120.690 131.125 120.860 ;
        RECT 131.720 120.590 132.120 121.190 ;
        RECT 128.605 120.440 128.775 120.475 ;
        RECT 128.520 119.590 128.870 120.440 ;
        RECT 128.520 119.190 129.520 119.590 ;
        RECT 129.895 119.435 130.065 120.475 ;
        RECT 131.185 120.440 131.355 120.475 ;
        RECT 131.120 119.590 131.420 120.440 ;
        RECT 129.220 118.790 129.520 119.190 ;
        RECT 130.420 119.190 131.420 119.590 ;
        RECT 131.720 119.290 133.120 120.590 ;
        RECT 130.420 118.790 130.720 119.190 ;
        RECT 129.220 118.390 130.720 118.790 ;
        RECT 127.870 116.290 128.220 118.190 ;
        RECT 128.520 117.190 128.870 118.190 ;
        RECT 128.605 116.955 128.775 117.190 ;
        RECT 129.720 116.990 130.220 118.390 ;
        RECT 131.120 117.190 131.420 118.190 ;
        RECT 129.895 116.955 130.065 116.990 ;
        RECT 131.185 116.955 131.355 117.190 ;
        RECT 131.720 116.890 133.120 118.190 ;
        RECT 128.835 116.615 129.835 116.785 ;
        RECT 130.125 116.615 131.125 116.785 ;
        RECT 131.720 116.290 132.120 116.890 ;
        RECT 127.870 115.940 132.120 116.290 ;
        RECT 127.010 113.365 132.070 113.535 ;
        RECT 127.265 112.565 127.520 113.365 ;
        RECT 127.690 112.395 128.020 113.195 ;
        RECT 128.190 112.565 128.360 113.365 ;
        RECT 128.530 112.395 128.860 113.195 ;
        RECT 129.030 112.565 129.200 113.365 ;
        RECT 129.370 112.395 129.700 113.195 ;
        RECT 129.870 112.565 130.040 113.365 ;
        RECT 130.210 112.395 130.540 113.195 ;
        RECT 130.710 112.565 131.010 113.365 ;
        RECT 127.095 112.225 131.065 112.395 ;
        RECT 127.095 111.635 127.440 112.225 ;
        RECT 127.690 111.805 130.545 112.055 ;
        RECT 130.745 111.635 131.065 112.225 ;
        RECT 131.235 112.200 131.985 113.185 ;
        RECT 127.095 111.445 131.065 111.635 ;
        RECT 127.265 110.815 127.520 111.275 ;
        RECT 127.690 110.985 128.020 111.445 ;
        RECT 128.190 110.815 128.360 111.275 ;
        RECT 128.530 110.985 128.860 111.445 ;
        RECT 129.030 110.815 129.200 111.275 ;
        RECT 129.370 110.985 129.700 111.445 ;
        RECT 129.870 110.815 130.040 111.275 ;
        RECT 130.210 110.985 130.540 111.445 ;
        RECT 130.710 110.815 131.015 111.275 ;
        RECT 131.235 110.995 131.985 111.540 ;
        RECT 127.010 110.645 132.070 110.815 ;
        RECT 111.700 109.490 123.550 109.640 ;
        RECT 111.700 109.470 121.160 109.490 ;
        RECT 121.900 109.470 123.550 109.490 ;
        RECT 63.710 93.910 67.960 94.160 ;
        RECT 63.710 91.910 64.060 93.910 ;
        RECT 64.675 93.410 65.675 93.580 ;
        RECT 65.965 93.410 66.965 93.580 ;
        RECT 67.560 93.310 67.960 93.910 ;
        RECT 64.445 93.160 64.615 93.195 ;
        RECT 64.360 92.310 64.710 93.160 ;
        RECT 64.360 91.910 65.360 92.310 ;
        RECT 65.735 92.155 65.905 93.195 ;
        RECT 67.025 93.160 67.195 93.195 ;
        RECT 66.960 92.310 67.260 93.160 ;
        RECT 65.060 91.510 65.360 91.910 ;
        RECT 66.260 91.910 67.260 92.310 ;
        RECT 67.560 92.010 68.960 93.310 ;
        RECT 129.620 93.260 133.870 93.510 ;
        RECT 66.260 91.510 66.560 91.910 ;
        RECT 28.580 91.030 56.300 91.360 ;
        RECT 65.060 91.110 66.560 91.510 ;
        RECT 129.620 91.260 129.970 93.260 ;
        RECT 130.585 92.760 131.585 92.930 ;
        RECT 131.875 92.760 132.875 92.930 ;
        RECT 133.470 92.660 133.870 93.260 ;
        RECT 130.355 92.510 130.525 92.545 ;
        RECT 130.270 91.660 130.620 92.510 ;
        RECT 130.270 91.260 131.270 91.660 ;
        RECT 131.645 91.505 131.815 92.545 ;
        RECT 132.935 92.510 133.105 92.545 ;
        RECT 132.870 91.660 133.170 92.510 ;
        RECT 28.580 78.160 28.910 91.030 ;
        RECT 29.900 89.380 54.980 89.710 ;
        RECT 29.900 79.810 30.230 89.380 ;
        RECT 34.760 87.410 53.210 88.010 ;
        RECT 37.530 86.150 37.700 87.190 ;
        RECT 38.820 86.150 38.990 87.190 ;
        RECT 40.110 86.150 40.280 87.190 ;
        RECT 41.400 86.150 41.570 87.190 ;
        RECT 42.690 86.150 42.860 87.190 ;
        RECT 43.980 86.150 44.150 87.190 ;
        RECT 45.270 86.150 45.440 87.190 ;
        RECT 46.560 86.150 46.730 87.190 ;
        RECT 47.850 86.150 48.020 87.190 ;
        RECT 49.140 86.150 49.310 87.190 ;
        RECT 50.430 86.150 50.600 87.190 ;
        RECT 51.720 86.150 51.890 87.190 ;
        RECT 53.010 86.150 53.180 87.190 ;
        RECT 37.760 85.765 38.760 85.935 ;
        RECT 39.050 85.765 40.050 85.935 ;
        RECT 40.340 85.765 41.340 85.935 ;
        RECT 41.630 85.765 42.630 85.935 ;
        RECT 42.920 85.765 43.920 85.935 ;
        RECT 44.210 85.765 45.210 85.935 ;
        RECT 45.500 85.765 46.500 85.935 ;
        RECT 46.790 85.765 47.790 85.935 ;
        RECT 48.080 85.765 49.080 85.935 ;
        RECT 49.370 85.765 50.370 85.935 ;
        RECT 50.660 85.765 51.660 85.935 ;
        RECT 51.950 85.765 52.950 85.935 ;
        RECT 39.050 85.225 40.050 85.395 ;
        RECT 42.920 85.225 43.920 85.395 ;
        RECT 44.210 85.225 45.210 85.395 ;
        RECT 48.080 85.225 49.080 85.395 ;
        RECT 49.370 85.225 50.370 85.395 ;
        RECT 37.530 84.015 37.700 85.055 ;
        RECT 38.820 84.015 38.990 85.055 ;
        RECT 40.110 84.015 40.280 85.055 ;
        RECT 41.400 84.015 41.570 85.055 ;
        RECT 42.690 84.015 42.860 85.055 ;
        RECT 43.980 84.015 44.150 85.055 ;
        RECT 45.270 84.015 45.440 85.055 ;
        RECT 46.560 84.015 46.730 85.055 ;
        RECT 47.850 84.015 48.020 85.055 ;
        RECT 49.140 84.015 49.310 85.055 ;
        RECT 50.430 84.015 50.600 85.055 ;
        RECT 51.720 84.015 51.890 85.055 ;
        RECT 53.010 84.015 53.180 85.055 ;
        RECT 37.760 83.675 38.760 83.845 ;
        RECT 40.340 83.675 41.340 83.845 ;
        RECT 41.630 83.675 42.630 83.845 ;
        RECT 45.500 83.675 46.500 83.845 ;
        RECT 46.790 83.675 47.790 83.845 ;
        RECT 50.660 83.675 51.660 83.845 ;
        RECT 51.950 83.675 52.950 83.845 ;
        RECT 37.760 83.045 38.760 83.215 ;
        RECT 39.050 83.045 40.050 83.215 ;
        RECT 40.340 83.045 41.340 83.215 ;
        RECT 41.630 83.045 42.630 83.215 ;
        RECT 42.920 83.045 43.920 83.215 ;
        RECT 44.210 83.045 45.210 83.215 ;
        RECT 45.500 83.045 46.500 83.215 ;
        RECT 46.790 83.045 47.790 83.215 ;
        RECT 48.080 83.045 49.080 83.215 ;
        RECT 49.370 83.045 50.370 83.215 ;
        RECT 50.660 83.045 51.660 83.215 ;
        RECT 51.950 83.045 52.950 83.215 ;
        RECT 37.530 82.415 37.700 82.875 ;
        RECT 38.820 82.415 38.990 82.875 ;
        RECT 40.110 82.415 40.280 82.875 ;
        RECT 41.400 82.415 41.570 82.875 ;
        RECT 42.690 82.415 42.860 82.875 ;
        RECT 43.980 82.415 44.150 82.875 ;
        RECT 45.270 82.415 45.440 82.875 ;
        RECT 46.560 82.415 46.730 82.875 ;
        RECT 47.850 82.415 48.020 82.875 ;
        RECT 49.140 82.415 49.310 82.875 ;
        RECT 50.430 82.415 50.600 82.875 ;
        RECT 51.720 82.415 51.890 82.875 ;
        RECT 53.010 82.415 53.180 82.875 ;
        RECT 34.760 81.610 36.960 82.310 ;
        RECT 37.510 81.460 53.210 82.010 ;
        RECT 54.650 79.810 54.980 89.380 ;
        RECT 29.900 79.480 54.980 79.810 ;
        RECT 55.970 78.160 56.300 91.030 ;
        RECT 57.740 90.180 59.390 90.350 ;
        RECT 57.740 82.010 57.910 90.180 ;
        RECT 58.160 87.510 58.960 89.710 ;
        RECT 57.160 79.610 57.910 82.010 ;
        RECT 28.580 77.830 56.300 78.160 ;
        RECT 47.660 76.540 53.460 77.010 ;
        RECT 47.540 76.510 57.000 76.540 ;
        RECT 57.740 76.510 57.910 79.610 ;
        RECT 47.540 76.370 57.910 76.510 ;
        RECT 47.540 75.060 47.710 76.370 ;
        RECT 48.190 75.540 50.350 75.890 ;
        RECT 54.190 75.540 56.350 75.890 ;
        RECT 56.830 75.060 57.910 76.370 ;
        RECT 58.390 75.540 58.740 77.700 ;
        RECT 59.220 75.060 59.390 90.180 ;
        RECT 63.710 89.010 64.060 90.910 ;
        RECT 64.360 89.910 64.710 90.910 ;
        RECT 64.445 89.675 64.615 89.910 ;
        RECT 65.560 89.710 66.060 91.110 ;
        RECT 66.960 89.910 67.260 90.910 ;
        RECT 65.735 89.675 65.905 89.710 ;
        RECT 67.025 89.675 67.195 89.910 ;
        RECT 67.560 89.610 68.960 90.910 ;
        RECT 130.970 90.860 131.270 91.260 ;
        RECT 132.170 91.260 133.170 91.660 ;
        RECT 133.470 91.360 134.870 92.660 ;
        RECT 132.170 90.860 132.470 91.260 ;
        RECT 94.490 90.380 122.210 90.710 ;
        RECT 130.970 90.460 132.470 90.860 ;
        RECT 64.675 89.335 65.675 89.505 ;
        RECT 65.965 89.335 66.965 89.505 ;
        RECT 67.560 89.010 67.960 89.610 ;
        RECT 63.710 88.660 67.960 89.010 ;
        RECT 63.710 86.610 67.960 86.860 ;
        RECT 63.710 84.610 64.060 86.610 ;
        RECT 64.675 86.110 65.675 86.280 ;
        RECT 65.965 86.110 66.965 86.280 ;
        RECT 67.560 86.010 67.960 86.610 ;
        RECT 64.445 85.860 64.615 85.895 ;
        RECT 64.360 85.010 64.710 85.860 ;
        RECT 64.360 84.610 65.360 85.010 ;
        RECT 65.735 84.855 65.905 85.895 ;
        RECT 67.025 85.860 67.195 85.895 ;
        RECT 66.960 85.010 67.260 85.860 ;
        RECT 65.060 84.210 65.360 84.610 ;
        RECT 66.260 84.610 67.260 85.010 ;
        RECT 67.560 84.710 68.960 86.010 ;
        RECT 66.260 84.210 66.560 84.610 ;
        RECT 65.060 83.810 66.560 84.210 ;
        RECT 63.710 81.710 64.060 83.610 ;
        RECT 64.360 82.610 64.710 83.610 ;
        RECT 64.445 82.375 64.615 82.610 ;
        RECT 65.560 82.410 66.060 83.810 ;
        RECT 66.960 82.610 67.260 83.610 ;
        RECT 65.735 82.375 65.905 82.410 ;
        RECT 67.025 82.375 67.195 82.610 ;
        RECT 67.560 82.310 68.960 83.610 ;
        RECT 64.675 82.035 65.675 82.205 ;
        RECT 65.965 82.035 66.965 82.205 ;
        RECT 67.560 81.710 67.960 82.310 ;
        RECT 63.710 81.360 67.960 81.710 ;
        RECT 62.850 78.785 67.910 78.955 ;
        RECT 63.105 77.985 63.360 78.785 ;
        RECT 63.530 77.815 63.860 78.615 ;
        RECT 64.030 77.985 64.200 78.785 ;
        RECT 64.370 77.815 64.700 78.615 ;
        RECT 64.870 77.985 65.040 78.785 ;
        RECT 65.210 77.815 65.540 78.615 ;
        RECT 65.710 77.985 65.880 78.785 ;
        RECT 66.050 77.815 66.380 78.615 ;
        RECT 66.550 77.985 66.850 78.785 ;
        RECT 62.935 77.645 66.905 77.815 ;
        RECT 62.935 77.055 63.280 77.645 ;
        RECT 63.530 77.225 66.385 77.475 ;
        RECT 66.585 77.055 66.905 77.645 ;
        RECT 67.075 77.620 67.825 78.605 ;
        RECT 94.490 77.510 94.820 90.380 ;
        RECT 95.810 88.730 120.890 89.060 ;
        RECT 95.810 79.160 96.140 88.730 ;
        RECT 100.670 86.760 119.120 87.360 ;
        RECT 103.440 85.500 103.610 86.540 ;
        RECT 104.730 85.500 104.900 86.540 ;
        RECT 106.020 85.500 106.190 86.540 ;
        RECT 107.310 85.500 107.480 86.540 ;
        RECT 108.600 85.500 108.770 86.540 ;
        RECT 109.890 85.500 110.060 86.540 ;
        RECT 111.180 85.500 111.350 86.540 ;
        RECT 112.470 85.500 112.640 86.540 ;
        RECT 113.760 85.500 113.930 86.540 ;
        RECT 115.050 85.500 115.220 86.540 ;
        RECT 116.340 85.500 116.510 86.540 ;
        RECT 117.630 85.500 117.800 86.540 ;
        RECT 118.920 85.500 119.090 86.540 ;
        RECT 103.670 85.115 104.670 85.285 ;
        RECT 104.960 85.115 105.960 85.285 ;
        RECT 106.250 85.115 107.250 85.285 ;
        RECT 107.540 85.115 108.540 85.285 ;
        RECT 108.830 85.115 109.830 85.285 ;
        RECT 110.120 85.115 111.120 85.285 ;
        RECT 111.410 85.115 112.410 85.285 ;
        RECT 112.700 85.115 113.700 85.285 ;
        RECT 113.990 85.115 114.990 85.285 ;
        RECT 115.280 85.115 116.280 85.285 ;
        RECT 116.570 85.115 117.570 85.285 ;
        RECT 117.860 85.115 118.860 85.285 ;
        RECT 104.960 84.575 105.960 84.745 ;
        RECT 108.830 84.575 109.830 84.745 ;
        RECT 110.120 84.575 111.120 84.745 ;
        RECT 113.990 84.575 114.990 84.745 ;
        RECT 115.280 84.575 116.280 84.745 ;
        RECT 103.440 83.365 103.610 84.405 ;
        RECT 104.730 83.365 104.900 84.405 ;
        RECT 106.020 83.365 106.190 84.405 ;
        RECT 107.310 83.365 107.480 84.405 ;
        RECT 108.600 83.365 108.770 84.405 ;
        RECT 109.890 83.365 110.060 84.405 ;
        RECT 111.180 83.365 111.350 84.405 ;
        RECT 112.470 83.365 112.640 84.405 ;
        RECT 113.760 83.365 113.930 84.405 ;
        RECT 115.050 83.365 115.220 84.405 ;
        RECT 116.340 83.365 116.510 84.405 ;
        RECT 117.630 83.365 117.800 84.405 ;
        RECT 118.920 83.365 119.090 84.405 ;
        RECT 103.670 83.025 104.670 83.195 ;
        RECT 106.250 83.025 107.250 83.195 ;
        RECT 107.540 83.025 108.540 83.195 ;
        RECT 111.410 83.025 112.410 83.195 ;
        RECT 112.700 83.025 113.700 83.195 ;
        RECT 116.570 83.025 117.570 83.195 ;
        RECT 117.860 83.025 118.860 83.195 ;
        RECT 103.670 82.395 104.670 82.565 ;
        RECT 104.960 82.395 105.960 82.565 ;
        RECT 106.250 82.395 107.250 82.565 ;
        RECT 107.540 82.395 108.540 82.565 ;
        RECT 108.830 82.395 109.830 82.565 ;
        RECT 110.120 82.395 111.120 82.565 ;
        RECT 111.410 82.395 112.410 82.565 ;
        RECT 112.700 82.395 113.700 82.565 ;
        RECT 113.990 82.395 114.990 82.565 ;
        RECT 115.280 82.395 116.280 82.565 ;
        RECT 116.570 82.395 117.570 82.565 ;
        RECT 117.860 82.395 118.860 82.565 ;
        RECT 103.440 81.765 103.610 82.225 ;
        RECT 104.730 81.765 104.900 82.225 ;
        RECT 106.020 81.765 106.190 82.225 ;
        RECT 107.310 81.765 107.480 82.225 ;
        RECT 108.600 81.765 108.770 82.225 ;
        RECT 109.890 81.765 110.060 82.225 ;
        RECT 111.180 81.765 111.350 82.225 ;
        RECT 112.470 81.765 112.640 82.225 ;
        RECT 113.760 81.765 113.930 82.225 ;
        RECT 115.050 81.765 115.220 82.225 ;
        RECT 116.340 81.765 116.510 82.225 ;
        RECT 117.630 81.765 117.800 82.225 ;
        RECT 118.920 81.765 119.090 82.225 ;
        RECT 100.670 80.960 102.870 81.660 ;
        RECT 103.420 80.810 119.120 81.360 ;
        RECT 120.560 79.160 120.890 88.730 ;
        RECT 95.810 78.830 120.890 79.160 ;
        RECT 121.880 77.510 122.210 90.380 ;
        RECT 123.650 89.530 125.300 89.700 ;
        RECT 123.650 81.360 123.820 89.530 ;
        RECT 124.070 86.860 124.870 89.060 ;
        RECT 123.070 78.960 123.820 81.360 ;
        RECT 94.490 77.180 122.210 77.510 ;
        RECT 62.935 76.865 66.905 77.055 ;
        RECT 63.105 76.235 63.360 76.695 ;
        RECT 63.530 76.405 63.860 76.865 ;
        RECT 64.030 76.235 64.200 76.695 ;
        RECT 64.370 76.405 64.700 76.865 ;
        RECT 64.870 76.235 65.040 76.695 ;
        RECT 65.210 76.405 65.540 76.865 ;
        RECT 65.710 76.235 65.880 76.695 ;
        RECT 66.050 76.405 66.380 76.865 ;
        RECT 66.550 76.235 66.855 76.695 ;
        RECT 67.075 76.415 67.825 76.960 ;
        RECT 62.850 76.065 67.910 76.235 ;
        RECT 113.570 75.890 119.370 76.360 ;
        RECT 47.540 74.910 59.390 75.060 ;
        RECT 47.540 74.890 57.000 74.910 ;
        RECT 57.740 74.890 59.390 74.910 ;
        RECT 113.450 75.860 122.910 75.890 ;
        RECT 123.650 75.860 123.820 78.960 ;
        RECT 113.450 75.720 123.820 75.860 ;
        RECT 113.450 74.410 113.620 75.720 ;
        RECT 114.100 74.890 116.260 75.240 ;
        RECT 120.100 74.890 122.260 75.240 ;
        RECT 122.740 74.410 123.820 75.720 ;
        RECT 124.300 74.890 124.650 77.050 ;
        RECT 125.130 74.410 125.300 89.530 ;
        RECT 129.620 88.360 129.970 90.260 ;
        RECT 130.270 89.260 130.620 90.260 ;
        RECT 130.355 89.025 130.525 89.260 ;
        RECT 131.470 89.060 131.970 90.460 ;
        RECT 132.870 89.260 133.170 90.260 ;
        RECT 131.645 89.025 131.815 89.060 ;
        RECT 132.935 89.025 133.105 89.260 ;
        RECT 133.470 88.960 134.870 90.260 ;
        RECT 130.585 88.685 131.585 88.855 ;
        RECT 131.875 88.685 132.875 88.855 ;
        RECT 133.470 88.360 133.870 88.960 ;
        RECT 129.620 88.010 133.870 88.360 ;
        RECT 129.620 85.960 133.870 86.210 ;
        RECT 129.620 83.960 129.970 85.960 ;
        RECT 130.585 85.460 131.585 85.630 ;
        RECT 131.875 85.460 132.875 85.630 ;
        RECT 133.470 85.360 133.870 85.960 ;
        RECT 130.355 85.210 130.525 85.245 ;
        RECT 130.270 84.360 130.620 85.210 ;
        RECT 130.270 83.960 131.270 84.360 ;
        RECT 131.645 84.205 131.815 85.245 ;
        RECT 132.935 85.210 133.105 85.245 ;
        RECT 132.870 84.360 133.170 85.210 ;
        RECT 130.970 83.560 131.270 83.960 ;
        RECT 132.170 83.960 133.170 84.360 ;
        RECT 133.470 84.060 134.870 85.360 ;
        RECT 132.170 83.560 132.470 83.960 ;
        RECT 130.970 83.160 132.470 83.560 ;
        RECT 129.620 81.060 129.970 82.960 ;
        RECT 130.270 81.960 130.620 82.960 ;
        RECT 130.355 81.725 130.525 81.960 ;
        RECT 131.470 81.760 131.970 83.160 ;
        RECT 132.870 81.960 133.170 82.960 ;
        RECT 131.645 81.725 131.815 81.760 ;
        RECT 132.935 81.725 133.105 81.960 ;
        RECT 133.470 81.660 134.870 82.960 ;
        RECT 130.585 81.385 131.585 81.555 ;
        RECT 131.875 81.385 132.875 81.555 ;
        RECT 133.470 81.060 133.870 81.660 ;
        RECT 129.620 80.710 133.870 81.060 ;
        RECT 128.760 78.135 133.820 78.305 ;
        RECT 129.015 77.335 129.270 78.135 ;
        RECT 129.440 77.165 129.770 77.965 ;
        RECT 129.940 77.335 130.110 78.135 ;
        RECT 130.280 77.165 130.610 77.965 ;
        RECT 130.780 77.335 130.950 78.135 ;
        RECT 131.120 77.165 131.450 77.965 ;
        RECT 131.620 77.335 131.790 78.135 ;
        RECT 131.960 77.165 132.290 77.965 ;
        RECT 132.460 77.335 132.760 78.135 ;
        RECT 128.845 76.995 132.815 77.165 ;
        RECT 128.845 76.405 129.190 76.995 ;
        RECT 129.440 76.575 132.295 76.825 ;
        RECT 132.495 76.405 132.815 76.995 ;
        RECT 132.985 76.970 133.735 77.955 ;
        RECT 128.845 76.215 132.815 76.405 ;
        RECT 129.015 75.585 129.270 76.045 ;
        RECT 129.440 75.755 129.770 76.215 ;
        RECT 129.940 75.585 130.110 76.045 ;
        RECT 130.280 75.755 130.610 76.215 ;
        RECT 130.780 75.585 130.950 76.045 ;
        RECT 131.120 75.755 131.450 76.215 ;
        RECT 131.620 75.585 131.790 76.045 ;
        RECT 131.960 75.755 132.290 76.215 ;
        RECT 132.460 75.585 132.765 76.045 ;
        RECT 132.985 75.765 133.735 76.310 ;
        RECT 128.760 75.415 133.820 75.585 ;
        RECT 113.450 74.260 125.300 74.410 ;
        RECT 113.450 74.240 122.910 74.260 ;
        RECT 123.650 74.240 125.300 74.260 ;
      LAYER mcon ;
        RECT 64.545 191.600 65.385 191.770 ;
        RECT 65.835 191.600 66.675 191.770 ;
        RECT 64.235 190.425 64.405 191.305 ;
        RECT 65.525 190.425 65.695 191.305 ;
        RECT 66.815 190.425 66.985 191.305 ;
        RECT 68.150 190.400 68.650 191.300 ;
        RECT 128.615 192.380 129.455 192.550 ;
        RECT 129.905 192.380 130.745 192.550 ;
        RECT 128.305 191.205 128.475 192.085 ;
        RECT 129.595 191.205 129.765 192.085 ;
        RECT 130.885 191.205 131.055 192.085 ;
        RECT 132.220 191.180 132.720 192.080 ;
        RECT 28.450 189.300 56.050 189.500 ;
        RECT 28.450 176.300 28.650 189.300 ;
        RECT 29.750 187.650 54.700 187.850 ;
        RECT 29.750 177.950 29.950 187.650 ;
        RECT 34.850 185.800 52.750 186.000 ;
        RECT 37.320 184.420 37.490 185.300 ;
        RECT 38.610 184.420 38.780 185.300 ;
        RECT 39.900 184.420 40.070 185.300 ;
        RECT 41.190 184.420 41.360 185.300 ;
        RECT 42.480 184.420 42.650 185.300 ;
        RECT 43.770 184.420 43.940 185.300 ;
        RECT 45.060 184.420 45.230 185.300 ;
        RECT 46.350 184.420 46.520 185.300 ;
        RECT 47.640 184.420 47.810 185.300 ;
        RECT 48.930 184.420 49.100 185.300 ;
        RECT 50.220 184.420 50.390 185.300 ;
        RECT 51.510 184.420 51.680 185.300 ;
        RECT 52.800 184.420 52.970 185.300 ;
        RECT 37.630 183.955 38.470 184.125 ;
        RECT 38.920 183.955 39.760 184.125 ;
        RECT 40.210 183.955 41.050 184.125 ;
        RECT 41.500 183.955 42.340 184.125 ;
        RECT 42.790 183.955 43.630 184.125 ;
        RECT 44.080 183.955 44.920 184.125 ;
        RECT 45.370 183.955 46.210 184.125 ;
        RECT 46.660 183.955 47.500 184.125 ;
        RECT 47.950 183.955 48.790 184.125 ;
        RECT 49.240 183.955 50.080 184.125 ;
        RECT 50.530 183.955 51.370 184.125 ;
        RECT 51.820 183.955 52.660 184.125 ;
        RECT 38.920 183.415 39.760 183.585 ;
        RECT 42.790 183.415 43.630 183.585 ;
        RECT 44.080 183.415 44.920 183.585 ;
        RECT 47.950 183.415 48.790 183.585 ;
        RECT 49.240 183.415 50.080 183.585 ;
        RECT 37.320 182.285 37.490 183.165 ;
        RECT 38.610 182.285 38.780 183.165 ;
        RECT 39.900 182.285 40.070 183.165 ;
        RECT 41.190 182.285 41.360 183.165 ;
        RECT 42.480 182.285 42.650 183.165 ;
        RECT 43.770 182.285 43.940 183.165 ;
        RECT 45.060 182.285 45.230 183.165 ;
        RECT 46.350 182.285 46.520 183.165 ;
        RECT 47.640 182.285 47.810 183.165 ;
        RECT 48.930 182.285 49.100 183.165 ;
        RECT 50.220 182.285 50.390 183.165 ;
        RECT 51.510 182.285 51.680 183.165 ;
        RECT 52.800 182.285 52.970 183.165 ;
        RECT 37.630 181.865 38.470 182.035 ;
        RECT 40.210 181.865 41.050 182.035 ;
        RECT 41.500 181.865 42.340 182.035 ;
        RECT 45.370 181.865 46.210 182.035 ;
        RECT 46.660 181.865 47.500 182.035 ;
        RECT 50.530 181.865 51.370 182.035 ;
        RECT 51.820 181.865 52.660 182.035 ;
        RECT 37.630 181.235 38.470 181.405 ;
        RECT 38.920 181.235 39.760 181.405 ;
        RECT 40.210 181.235 41.050 181.405 ;
        RECT 41.500 181.235 42.340 181.405 ;
        RECT 42.790 181.235 43.630 181.405 ;
        RECT 44.080 181.235 44.920 181.405 ;
        RECT 45.370 181.235 46.210 181.405 ;
        RECT 46.660 181.235 47.500 181.405 ;
        RECT 47.950 181.235 48.790 181.405 ;
        RECT 49.240 181.235 50.080 181.405 ;
        RECT 50.530 181.235 51.370 181.405 ;
        RECT 51.820 181.235 52.660 181.405 ;
        RECT 37.320 180.685 37.490 180.985 ;
        RECT 38.610 180.685 38.780 180.985 ;
        RECT 39.900 180.685 40.070 180.985 ;
        RECT 41.190 180.685 41.360 180.985 ;
        RECT 42.480 180.685 42.650 180.985 ;
        RECT 43.770 180.685 43.940 180.985 ;
        RECT 45.060 180.685 45.230 180.985 ;
        RECT 46.350 180.685 46.520 180.985 ;
        RECT 47.640 180.685 47.810 180.985 ;
        RECT 48.930 180.685 49.100 180.985 ;
        RECT 50.220 180.685 50.390 180.985 ;
        RECT 51.510 180.685 51.680 180.985 ;
        RECT 52.800 180.685 52.970 180.985 ;
        RECT 34.650 179.900 36.650 180.350 ;
        RECT 37.500 179.800 52.750 180.050 ;
        RECT 54.500 177.950 54.700 187.650 ;
        RECT 29.750 177.750 54.700 177.950 ;
        RECT 55.850 176.300 56.050 189.300 ;
        RECT 28.450 176.100 56.050 176.300 ;
        RECT 58.050 185.800 58.650 187.800 ;
        RECT 57.050 177.900 57.550 180.100 ;
        RECT 47.550 174.700 53.150 175.100 ;
        RECT 48.070 173.810 50.055 174.000 ;
        RECT 54.065 173.810 56.050 174.000 ;
        RECT 58.260 173.820 58.450 175.805 ;
        RECT 64.235 187.945 64.405 188.825 ;
        RECT 65.525 187.945 65.695 188.825 ;
        RECT 66.815 187.945 66.985 188.825 ;
        RECT 68.150 188.000 68.650 188.900 ;
        RECT 64.545 187.525 65.385 187.695 ;
        RECT 65.835 187.525 66.675 187.695 ;
        RECT 64.545 184.300 65.385 184.470 ;
        RECT 65.835 184.300 66.675 184.470 ;
        RECT 64.235 183.125 64.405 184.005 ;
        RECT 65.525 183.125 65.695 184.005 ;
        RECT 66.815 183.125 66.985 184.005 ;
        RECT 68.150 183.100 68.650 184.000 ;
        RECT 64.235 180.645 64.405 181.525 ;
        RECT 65.525 180.645 65.695 181.525 ;
        RECT 66.815 180.645 66.985 181.525 ;
        RECT 68.150 180.700 68.650 181.600 ;
        RECT 64.545 180.225 65.385 180.395 ;
        RECT 65.835 180.225 66.675 180.395 ;
        RECT 62.785 176.975 62.955 177.145 ;
        RECT 63.245 176.975 63.415 177.145 ;
        RECT 63.705 176.975 63.875 177.145 ;
        RECT 64.165 176.975 64.335 177.145 ;
        RECT 64.625 176.975 64.795 177.145 ;
        RECT 65.085 176.975 65.255 177.145 ;
        RECT 65.545 176.975 65.715 177.145 ;
        RECT 66.005 176.975 66.175 177.145 ;
        RECT 66.465 176.975 66.635 177.145 ;
        RECT 66.925 176.975 67.095 177.145 ;
        RECT 67.385 176.975 67.555 177.145 ;
        RECT 92.520 190.080 120.120 190.280 ;
        RECT 92.520 177.080 92.720 190.080 ;
        RECT 93.820 188.430 118.770 188.630 ;
        RECT 93.820 178.730 94.020 188.430 ;
        RECT 98.920 186.580 116.820 186.780 ;
        RECT 101.390 185.200 101.560 186.080 ;
        RECT 102.680 185.200 102.850 186.080 ;
        RECT 103.970 185.200 104.140 186.080 ;
        RECT 105.260 185.200 105.430 186.080 ;
        RECT 106.550 185.200 106.720 186.080 ;
        RECT 107.840 185.200 108.010 186.080 ;
        RECT 109.130 185.200 109.300 186.080 ;
        RECT 110.420 185.200 110.590 186.080 ;
        RECT 111.710 185.200 111.880 186.080 ;
        RECT 113.000 185.200 113.170 186.080 ;
        RECT 114.290 185.200 114.460 186.080 ;
        RECT 115.580 185.200 115.750 186.080 ;
        RECT 116.870 185.200 117.040 186.080 ;
        RECT 101.700 184.735 102.540 184.905 ;
        RECT 102.990 184.735 103.830 184.905 ;
        RECT 104.280 184.735 105.120 184.905 ;
        RECT 105.570 184.735 106.410 184.905 ;
        RECT 106.860 184.735 107.700 184.905 ;
        RECT 108.150 184.735 108.990 184.905 ;
        RECT 109.440 184.735 110.280 184.905 ;
        RECT 110.730 184.735 111.570 184.905 ;
        RECT 112.020 184.735 112.860 184.905 ;
        RECT 113.310 184.735 114.150 184.905 ;
        RECT 114.600 184.735 115.440 184.905 ;
        RECT 115.890 184.735 116.730 184.905 ;
        RECT 102.990 184.195 103.830 184.365 ;
        RECT 106.860 184.195 107.700 184.365 ;
        RECT 108.150 184.195 108.990 184.365 ;
        RECT 112.020 184.195 112.860 184.365 ;
        RECT 113.310 184.195 114.150 184.365 ;
        RECT 101.390 183.065 101.560 183.945 ;
        RECT 102.680 183.065 102.850 183.945 ;
        RECT 103.970 183.065 104.140 183.945 ;
        RECT 105.260 183.065 105.430 183.945 ;
        RECT 106.550 183.065 106.720 183.945 ;
        RECT 107.840 183.065 108.010 183.945 ;
        RECT 109.130 183.065 109.300 183.945 ;
        RECT 110.420 183.065 110.590 183.945 ;
        RECT 111.710 183.065 111.880 183.945 ;
        RECT 113.000 183.065 113.170 183.945 ;
        RECT 114.290 183.065 114.460 183.945 ;
        RECT 115.580 183.065 115.750 183.945 ;
        RECT 116.870 183.065 117.040 183.945 ;
        RECT 101.700 182.645 102.540 182.815 ;
        RECT 104.280 182.645 105.120 182.815 ;
        RECT 105.570 182.645 106.410 182.815 ;
        RECT 109.440 182.645 110.280 182.815 ;
        RECT 110.730 182.645 111.570 182.815 ;
        RECT 114.600 182.645 115.440 182.815 ;
        RECT 115.890 182.645 116.730 182.815 ;
        RECT 101.700 182.015 102.540 182.185 ;
        RECT 102.990 182.015 103.830 182.185 ;
        RECT 104.280 182.015 105.120 182.185 ;
        RECT 105.570 182.015 106.410 182.185 ;
        RECT 106.860 182.015 107.700 182.185 ;
        RECT 108.150 182.015 108.990 182.185 ;
        RECT 109.440 182.015 110.280 182.185 ;
        RECT 110.730 182.015 111.570 182.185 ;
        RECT 112.020 182.015 112.860 182.185 ;
        RECT 113.310 182.015 114.150 182.185 ;
        RECT 114.600 182.015 115.440 182.185 ;
        RECT 115.890 182.015 116.730 182.185 ;
        RECT 101.390 181.465 101.560 181.765 ;
        RECT 102.680 181.465 102.850 181.765 ;
        RECT 103.970 181.465 104.140 181.765 ;
        RECT 105.260 181.465 105.430 181.765 ;
        RECT 106.550 181.465 106.720 181.765 ;
        RECT 107.840 181.465 108.010 181.765 ;
        RECT 109.130 181.465 109.300 181.765 ;
        RECT 110.420 181.465 110.590 181.765 ;
        RECT 111.710 181.465 111.880 181.765 ;
        RECT 113.000 181.465 113.170 181.765 ;
        RECT 114.290 181.465 114.460 181.765 ;
        RECT 115.580 181.465 115.750 181.765 ;
        RECT 116.870 181.465 117.040 181.765 ;
        RECT 98.720 180.680 100.720 181.130 ;
        RECT 101.570 180.580 116.820 180.830 ;
        RECT 118.570 178.730 118.770 188.430 ;
        RECT 93.820 178.530 118.770 178.730 ;
        RECT 119.920 177.080 120.120 190.080 ;
        RECT 92.520 176.880 120.120 177.080 ;
        RECT 122.120 186.580 122.720 188.580 ;
        RECT 121.120 178.680 121.620 180.880 ;
        RECT 63.360 175.450 65.800 175.620 ;
        RECT 66.420 175.120 66.660 175.940 ;
        RECT 111.620 175.480 117.220 175.880 ;
        RECT 62.785 174.255 62.955 174.425 ;
        RECT 63.245 174.255 63.415 174.425 ;
        RECT 63.705 174.255 63.875 174.425 ;
        RECT 64.165 174.255 64.335 174.425 ;
        RECT 64.625 174.255 64.795 174.425 ;
        RECT 65.085 174.255 65.255 174.425 ;
        RECT 65.545 174.255 65.715 174.425 ;
        RECT 66.005 174.255 66.175 174.425 ;
        RECT 66.465 174.255 66.635 174.425 ;
        RECT 66.925 174.255 67.095 174.425 ;
        RECT 67.385 174.255 67.555 174.425 ;
        RECT 112.140 174.590 114.125 174.780 ;
        RECT 118.135 174.590 120.120 174.780 ;
        RECT 122.330 174.600 122.520 176.585 ;
        RECT 128.305 188.725 128.475 189.605 ;
        RECT 129.595 188.725 129.765 189.605 ;
        RECT 130.885 188.725 131.055 189.605 ;
        RECT 132.220 188.780 132.720 189.680 ;
        RECT 128.615 188.305 129.455 188.475 ;
        RECT 129.905 188.305 130.745 188.475 ;
        RECT 128.615 185.080 129.455 185.250 ;
        RECT 129.905 185.080 130.745 185.250 ;
        RECT 128.305 183.905 128.475 184.785 ;
        RECT 129.595 183.905 129.765 184.785 ;
        RECT 130.885 183.905 131.055 184.785 ;
        RECT 132.220 183.880 132.720 184.780 ;
        RECT 128.305 181.425 128.475 182.305 ;
        RECT 129.595 181.425 129.765 182.305 ;
        RECT 130.885 181.425 131.055 182.305 ;
        RECT 132.220 181.480 132.720 182.380 ;
        RECT 128.615 181.005 129.455 181.175 ;
        RECT 129.905 181.005 130.745 181.175 ;
        RECT 126.855 177.755 127.025 177.925 ;
        RECT 127.315 177.755 127.485 177.925 ;
        RECT 127.775 177.755 127.945 177.925 ;
        RECT 128.235 177.755 128.405 177.925 ;
        RECT 128.695 177.755 128.865 177.925 ;
        RECT 129.155 177.755 129.325 177.925 ;
        RECT 129.615 177.755 129.785 177.925 ;
        RECT 130.075 177.755 130.245 177.925 ;
        RECT 130.535 177.755 130.705 177.925 ;
        RECT 130.995 177.755 131.165 177.925 ;
        RECT 131.455 177.755 131.625 177.925 ;
        RECT 127.430 176.230 129.870 176.400 ;
        RECT 130.490 175.900 130.730 176.720 ;
        RECT 126.855 175.035 127.025 175.205 ;
        RECT 127.315 175.035 127.485 175.205 ;
        RECT 127.775 175.035 127.945 175.205 ;
        RECT 128.235 175.035 128.405 175.205 ;
        RECT 128.695 175.035 128.865 175.205 ;
        RECT 129.155 175.035 129.325 175.205 ;
        RECT 129.615 175.035 129.785 175.205 ;
        RECT 130.075 175.035 130.245 175.205 ;
        RECT 130.535 175.035 130.705 175.205 ;
        RECT 130.995 175.035 131.165 175.205 ;
        RECT 131.455 175.035 131.625 175.205 ;
        RECT 64.775 162.160 65.615 162.330 ;
        RECT 66.065 162.160 66.905 162.330 ;
        RECT 64.465 160.985 64.635 161.865 ;
        RECT 65.755 160.985 65.925 161.865 ;
        RECT 67.045 160.985 67.215 161.865 ;
        RECT 68.380 160.960 68.880 161.860 ;
        RECT 128.435 161.780 129.275 161.950 ;
        RECT 129.725 161.780 130.565 161.950 ;
        RECT 128.125 160.605 128.295 161.485 ;
        RECT 129.415 160.605 129.585 161.485 ;
        RECT 130.705 160.605 130.875 161.485 ;
        RECT 28.680 159.860 56.280 160.060 ;
        RECT 28.680 146.860 28.880 159.860 ;
        RECT 29.980 158.210 54.930 158.410 ;
        RECT 29.980 148.510 30.180 158.210 ;
        RECT 35.080 156.360 52.980 156.560 ;
        RECT 37.550 154.980 37.720 155.860 ;
        RECT 38.840 154.980 39.010 155.860 ;
        RECT 40.130 154.980 40.300 155.860 ;
        RECT 41.420 154.980 41.590 155.860 ;
        RECT 42.710 154.980 42.880 155.860 ;
        RECT 44.000 154.980 44.170 155.860 ;
        RECT 45.290 154.980 45.460 155.860 ;
        RECT 46.580 154.980 46.750 155.860 ;
        RECT 47.870 154.980 48.040 155.860 ;
        RECT 49.160 154.980 49.330 155.860 ;
        RECT 50.450 154.980 50.620 155.860 ;
        RECT 51.740 154.980 51.910 155.860 ;
        RECT 53.030 154.980 53.200 155.860 ;
        RECT 37.860 154.515 38.700 154.685 ;
        RECT 39.150 154.515 39.990 154.685 ;
        RECT 40.440 154.515 41.280 154.685 ;
        RECT 41.730 154.515 42.570 154.685 ;
        RECT 43.020 154.515 43.860 154.685 ;
        RECT 44.310 154.515 45.150 154.685 ;
        RECT 45.600 154.515 46.440 154.685 ;
        RECT 46.890 154.515 47.730 154.685 ;
        RECT 48.180 154.515 49.020 154.685 ;
        RECT 49.470 154.515 50.310 154.685 ;
        RECT 50.760 154.515 51.600 154.685 ;
        RECT 52.050 154.515 52.890 154.685 ;
        RECT 39.150 153.975 39.990 154.145 ;
        RECT 43.020 153.975 43.860 154.145 ;
        RECT 44.310 153.975 45.150 154.145 ;
        RECT 48.180 153.975 49.020 154.145 ;
        RECT 49.470 153.975 50.310 154.145 ;
        RECT 37.550 152.845 37.720 153.725 ;
        RECT 38.840 152.845 39.010 153.725 ;
        RECT 40.130 152.845 40.300 153.725 ;
        RECT 41.420 152.845 41.590 153.725 ;
        RECT 42.710 152.845 42.880 153.725 ;
        RECT 44.000 152.845 44.170 153.725 ;
        RECT 45.290 152.845 45.460 153.725 ;
        RECT 46.580 152.845 46.750 153.725 ;
        RECT 47.870 152.845 48.040 153.725 ;
        RECT 49.160 152.845 49.330 153.725 ;
        RECT 50.450 152.845 50.620 153.725 ;
        RECT 51.740 152.845 51.910 153.725 ;
        RECT 53.030 152.845 53.200 153.725 ;
        RECT 37.860 152.425 38.700 152.595 ;
        RECT 40.440 152.425 41.280 152.595 ;
        RECT 41.730 152.425 42.570 152.595 ;
        RECT 45.600 152.425 46.440 152.595 ;
        RECT 46.890 152.425 47.730 152.595 ;
        RECT 50.760 152.425 51.600 152.595 ;
        RECT 52.050 152.425 52.890 152.595 ;
        RECT 37.860 151.795 38.700 151.965 ;
        RECT 39.150 151.795 39.990 151.965 ;
        RECT 40.440 151.795 41.280 151.965 ;
        RECT 41.730 151.795 42.570 151.965 ;
        RECT 43.020 151.795 43.860 151.965 ;
        RECT 44.310 151.795 45.150 151.965 ;
        RECT 45.600 151.795 46.440 151.965 ;
        RECT 46.890 151.795 47.730 151.965 ;
        RECT 48.180 151.795 49.020 151.965 ;
        RECT 49.470 151.795 50.310 151.965 ;
        RECT 50.760 151.795 51.600 151.965 ;
        RECT 52.050 151.795 52.890 151.965 ;
        RECT 37.550 151.245 37.720 151.545 ;
        RECT 38.840 151.245 39.010 151.545 ;
        RECT 40.130 151.245 40.300 151.545 ;
        RECT 41.420 151.245 41.590 151.545 ;
        RECT 42.710 151.245 42.880 151.545 ;
        RECT 44.000 151.245 44.170 151.545 ;
        RECT 45.290 151.245 45.460 151.545 ;
        RECT 46.580 151.245 46.750 151.545 ;
        RECT 47.870 151.245 48.040 151.545 ;
        RECT 49.160 151.245 49.330 151.545 ;
        RECT 50.450 151.245 50.620 151.545 ;
        RECT 51.740 151.245 51.910 151.545 ;
        RECT 53.030 151.245 53.200 151.545 ;
        RECT 34.880 150.460 36.880 150.910 ;
        RECT 37.730 150.360 52.980 150.610 ;
        RECT 54.730 148.510 54.930 158.210 ;
        RECT 29.980 148.310 54.930 148.510 ;
        RECT 56.080 146.860 56.280 159.860 ;
        RECT 28.680 146.660 56.280 146.860 ;
        RECT 132.040 160.580 132.540 161.480 ;
        RECT 58.280 156.360 58.880 158.360 ;
        RECT 57.280 148.460 57.780 150.660 ;
        RECT 47.780 145.260 53.380 145.660 ;
        RECT 48.300 144.370 50.285 144.560 ;
        RECT 54.295 144.370 56.280 144.560 ;
        RECT 58.490 144.380 58.680 146.365 ;
        RECT 64.465 158.505 64.635 159.385 ;
        RECT 65.755 158.505 65.925 159.385 ;
        RECT 67.045 158.505 67.215 159.385 ;
        RECT 68.380 158.560 68.880 159.460 ;
        RECT 64.775 158.085 65.615 158.255 ;
        RECT 66.065 158.085 66.905 158.255 ;
        RECT 64.775 154.860 65.615 155.030 ;
        RECT 66.065 154.860 66.905 155.030 ;
        RECT 64.465 153.685 64.635 154.565 ;
        RECT 65.755 153.685 65.925 154.565 ;
        RECT 67.045 153.685 67.215 154.565 ;
        RECT 68.380 153.660 68.880 154.560 ;
        RECT 64.465 151.205 64.635 152.085 ;
        RECT 65.755 151.205 65.925 152.085 ;
        RECT 67.045 151.205 67.215 152.085 ;
        RECT 68.380 151.260 68.880 152.160 ;
        RECT 64.775 150.785 65.615 150.955 ;
        RECT 66.065 150.785 66.905 150.955 ;
        RECT 63.015 147.535 63.185 147.705 ;
        RECT 63.475 147.535 63.645 147.705 ;
        RECT 63.935 147.535 64.105 147.705 ;
        RECT 64.395 147.535 64.565 147.705 ;
        RECT 64.855 147.535 65.025 147.705 ;
        RECT 65.315 147.535 65.485 147.705 ;
        RECT 65.775 147.535 65.945 147.705 ;
        RECT 66.235 147.535 66.405 147.705 ;
        RECT 66.695 147.535 66.865 147.705 ;
        RECT 67.155 147.535 67.325 147.705 ;
        RECT 67.615 147.535 67.785 147.705 ;
        RECT 63.590 146.010 66.030 146.180 ;
        RECT 66.650 145.680 66.890 146.500 ;
        RECT 92.340 159.480 119.940 159.680 ;
        RECT 92.340 146.480 92.540 159.480 ;
        RECT 93.640 157.830 118.590 158.030 ;
        RECT 93.640 148.130 93.840 157.830 ;
        RECT 98.740 155.980 116.640 156.180 ;
        RECT 101.210 154.600 101.380 155.480 ;
        RECT 102.500 154.600 102.670 155.480 ;
        RECT 103.790 154.600 103.960 155.480 ;
        RECT 105.080 154.600 105.250 155.480 ;
        RECT 106.370 154.600 106.540 155.480 ;
        RECT 107.660 154.600 107.830 155.480 ;
        RECT 108.950 154.600 109.120 155.480 ;
        RECT 110.240 154.600 110.410 155.480 ;
        RECT 111.530 154.600 111.700 155.480 ;
        RECT 112.820 154.600 112.990 155.480 ;
        RECT 114.110 154.600 114.280 155.480 ;
        RECT 115.400 154.600 115.570 155.480 ;
        RECT 116.690 154.600 116.860 155.480 ;
        RECT 101.520 154.135 102.360 154.305 ;
        RECT 102.810 154.135 103.650 154.305 ;
        RECT 104.100 154.135 104.940 154.305 ;
        RECT 105.390 154.135 106.230 154.305 ;
        RECT 106.680 154.135 107.520 154.305 ;
        RECT 107.970 154.135 108.810 154.305 ;
        RECT 109.260 154.135 110.100 154.305 ;
        RECT 110.550 154.135 111.390 154.305 ;
        RECT 111.840 154.135 112.680 154.305 ;
        RECT 113.130 154.135 113.970 154.305 ;
        RECT 114.420 154.135 115.260 154.305 ;
        RECT 115.710 154.135 116.550 154.305 ;
        RECT 102.810 153.595 103.650 153.765 ;
        RECT 106.680 153.595 107.520 153.765 ;
        RECT 107.970 153.595 108.810 153.765 ;
        RECT 111.840 153.595 112.680 153.765 ;
        RECT 113.130 153.595 113.970 153.765 ;
        RECT 101.210 152.465 101.380 153.345 ;
        RECT 102.500 152.465 102.670 153.345 ;
        RECT 103.790 152.465 103.960 153.345 ;
        RECT 105.080 152.465 105.250 153.345 ;
        RECT 106.370 152.465 106.540 153.345 ;
        RECT 107.660 152.465 107.830 153.345 ;
        RECT 108.950 152.465 109.120 153.345 ;
        RECT 110.240 152.465 110.410 153.345 ;
        RECT 111.530 152.465 111.700 153.345 ;
        RECT 112.820 152.465 112.990 153.345 ;
        RECT 114.110 152.465 114.280 153.345 ;
        RECT 115.400 152.465 115.570 153.345 ;
        RECT 116.690 152.465 116.860 153.345 ;
        RECT 101.520 152.045 102.360 152.215 ;
        RECT 104.100 152.045 104.940 152.215 ;
        RECT 105.390 152.045 106.230 152.215 ;
        RECT 109.260 152.045 110.100 152.215 ;
        RECT 110.550 152.045 111.390 152.215 ;
        RECT 114.420 152.045 115.260 152.215 ;
        RECT 115.710 152.045 116.550 152.215 ;
        RECT 101.520 151.415 102.360 151.585 ;
        RECT 102.810 151.415 103.650 151.585 ;
        RECT 104.100 151.415 104.940 151.585 ;
        RECT 105.390 151.415 106.230 151.585 ;
        RECT 106.680 151.415 107.520 151.585 ;
        RECT 107.970 151.415 108.810 151.585 ;
        RECT 109.260 151.415 110.100 151.585 ;
        RECT 110.550 151.415 111.390 151.585 ;
        RECT 111.840 151.415 112.680 151.585 ;
        RECT 113.130 151.415 113.970 151.585 ;
        RECT 114.420 151.415 115.260 151.585 ;
        RECT 115.710 151.415 116.550 151.585 ;
        RECT 101.210 150.865 101.380 151.165 ;
        RECT 102.500 150.865 102.670 151.165 ;
        RECT 103.790 150.865 103.960 151.165 ;
        RECT 105.080 150.865 105.250 151.165 ;
        RECT 106.370 150.865 106.540 151.165 ;
        RECT 107.660 150.865 107.830 151.165 ;
        RECT 108.950 150.865 109.120 151.165 ;
        RECT 110.240 150.865 110.410 151.165 ;
        RECT 111.530 150.865 111.700 151.165 ;
        RECT 112.820 150.865 112.990 151.165 ;
        RECT 114.110 150.865 114.280 151.165 ;
        RECT 115.400 150.865 115.570 151.165 ;
        RECT 116.690 150.865 116.860 151.165 ;
        RECT 98.540 150.080 100.540 150.530 ;
        RECT 101.390 149.980 116.640 150.230 ;
        RECT 118.390 148.130 118.590 157.830 ;
        RECT 93.640 147.930 118.590 148.130 ;
        RECT 119.740 146.480 119.940 159.480 ;
        RECT 92.340 146.280 119.940 146.480 ;
        RECT 121.940 155.980 122.540 157.980 ;
        RECT 120.940 148.080 121.440 150.280 ;
        RECT 63.015 144.815 63.185 144.985 ;
        RECT 63.475 144.815 63.645 144.985 ;
        RECT 63.935 144.815 64.105 144.985 ;
        RECT 64.395 144.815 64.565 144.985 ;
        RECT 64.855 144.815 65.025 144.985 ;
        RECT 65.315 144.815 65.485 144.985 ;
        RECT 65.775 144.815 65.945 144.985 ;
        RECT 66.235 144.815 66.405 144.985 ;
        RECT 66.695 144.815 66.865 144.985 ;
        RECT 67.155 144.815 67.325 144.985 ;
        RECT 67.615 144.815 67.785 144.985 ;
        RECT 111.440 144.880 117.040 145.280 ;
        RECT 111.960 143.990 113.945 144.180 ;
        RECT 117.955 143.990 119.940 144.180 ;
        RECT 122.150 144.000 122.340 145.985 ;
        RECT 128.125 158.125 128.295 159.005 ;
        RECT 129.415 158.125 129.585 159.005 ;
        RECT 130.705 158.125 130.875 159.005 ;
        RECT 132.040 158.180 132.540 159.080 ;
        RECT 128.435 157.705 129.275 157.875 ;
        RECT 129.725 157.705 130.565 157.875 ;
        RECT 128.435 154.480 129.275 154.650 ;
        RECT 129.725 154.480 130.565 154.650 ;
        RECT 128.125 153.305 128.295 154.185 ;
        RECT 129.415 153.305 129.585 154.185 ;
        RECT 130.705 153.305 130.875 154.185 ;
        RECT 132.040 153.280 132.540 154.180 ;
        RECT 128.125 150.825 128.295 151.705 ;
        RECT 129.415 150.825 129.585 151.705 ;
        RECT 130.705 150.825 130.875 151.705 ;
        RECT 132.040 150.880 132.540 151.780 ;
        RECT 128.435 150.405 129.275 150.575 ;
        RECT 129.725 150.405 130.565 150.575 ;
        RECT 126.675 147.155 126.845 147.325 ;
        RECT 127.135 147.155 127.305 147.325 ;
        RECT 127.595 147.155 127.765 147.325 ;
        RECT 128.055 147.155 128.225 147.325 ;
        RECT 128.515 147.155 128.685 147.325 ;
        RECT 128.975 147.155 129.145 147.325 ;
        RECT 129.435 147.155 129.605 147.325 ;
        RECT 129.895 147.155 130.065 147.325 ;
        RECT 130.355 147.155 130.525 147.325 ;
        RECT 130.815 147.155 130.985 147.325 ;
        RECT 131.275 147.155 131.445 147.325 ;
        RECT 127.250 145.630 129.690 145.800 ;
        RECT 130.310 145.300 130.550 146.120 ;
        RECT 126.675 144.435 126.845 144.605 ;
        RECT 127.135 144.435 127.305 144.605 ;
        RECT 127.595 144.435 127.765 144.605 ;
        RECT 128.055 144.435 128.225 144.605 ;
        RECT 128.515 144.435 128.685 144.605 ;
        RECT 128.975 144.435 129.145 144.605 ;
        RECT 129.435 144.435 129.605 144.605 ;
        RECT 129.895 144.435 130.065 144.605 ;
        RECT 130.355 144.435 130.525 144.605 ;
        RECT 130.815 144.435 130.985 144.605 ;
        RECT 131.275 144.435 131.445 144.605 ;
        RECT 65.375 128.640 66.215 128.810 ;
        RECT 66.665 128.640 67.505 128.810 ;
        RECT 65.065 127.465 65.235 128.345 ;
        RECT 66.355 127.465 66.525 128.345 ;
        RECT 67.645 127.465 67.815 128.345 ;
        RECT 68.980 127.440 69.480 128.340 ;
        RECT 29.280 126.340 56.880 126.540 ;
        RECT 29.280 113.340 29.480 126.340 ;
        RECT 30.580 124.690 55.530 124.890 ;
        RECT 30.580 114.990 30.780 124.690 ;
        RECT 35.680 122.840 53.580 123.040 ;
        RECT 38.150 121.460 38.320 122.340 ;
        RECT 39.440 121.460 39.610 122.340 ;
        RECT 40.730 121.460 40.900 122.340 ;
        RECT 42.020 121.460 42.190 122.340 ;
        RECT 43.310 121.460 43.480 122.340 ;
        RECT 44.600 121.460 44.770 122.340 ;
        RECT 45.890 121.460 46.060 122.340 ;
        RECT 47.180 121.460 47.350 122.340 ;
        RECT 48.470 121.460 48.640 122.340 ;
        RECT 49.760 121.460 49.930 122.340 ;
        RECT 51.050 121.460 51.220 122.340 ;
        RECT 52.340 121.460 52.510 122.340 ;
        RECT 53.630 121.460 53.800 122.340 ;
        RECT 38.460 120.995 39.300 121.165 ;
        RECT 39.750 120.995 40.590 121.165 ;
        RECT 41.040 120.995 41.880 121.165 ;
        RECT 42.330 120.995 43.170 121.165 ;
        RECT 43.620 120.995 44.460 121.165 ;
        RECT 44.910 120.995 45.750 121.165 ;
        RECT 46.200 120.995 47.040 121.165 ;
        RECT 47.490 120.995 48.330 121.165 ;
        RECT 48.780 120.995 49.620 121.165 ;
        RECT 50.070 120.995 50.910 121.165 ;
        RECT 51.360 120.995 52.200 121.165 ;
        RECT 52.650 120.995 53.490 121.165 ;
        RECT 39.750 120.455 40.590 120.625 ;
        RECT 43.620 120.455 44.460 120.625 ;
        RECT 44.910 120.455 45.750 120.625 ;
        RECT 48.780 120.455 49.620 120.625 ;
        RECT 50.070 120.455 50.910 120.625 ;
        RECT 38.150 119.325 38.320 120.205 ;
        RECT 39.440 119.325 39.610 120.205 ;
        RECT 40.730 119.325 40.900 120.205 ;
        RECT 42.020 119.325 42.190 120.205 ;
        RECT 43.310 119.325 43.480 120.205 ;
        RECT 44.600 119.325 44.770 120.205 ;
        RECT 45.890 119.325 46.060 120.205 ;
        RECT 47.180 119.325 47.350 120.205 ;
        RECT 48.470 119.325 48.640 120.205 ;
        RECT 49.760 119.325 49.930 120.205 ;
        RECT 51.050 119.325 51.220 120.205 ;
        RECT 52.340 119.325 52.510 120.205 ;
        RECT 53.630 119.325 53.800 120.205 ;
        RECT 38.460 118.905 39.300 119.075 ;
        RECT 41.040 118.905 41.880 119.075 ;
        RECT 42.330 118.905 43.170 119.075 ;
        RECT 46.200 118.905 47.040 119.075 ;
        RECT 47.490 118.905 48.330 119.075 ;
        RECT 51.360 118.905 52.200 119.075 ;
        RECT 52.650 118.905 53.490 119.075 ;
        RECT 38.460 118.275 39.300 118.445 ;
        RECT 39.750 118.275 40.590 118.445 ;
        RECT 41.040 118.275 41.880 118.445 ;
        RECT 42.330 118.275 43.170 118.445 ;
        RECT 43.620 118.275 44.460 118.445 ;
        RECT 44.910 118.275 45.750 118.445 ;
        RECT 46.200 118.275 47.040 118.445 ;
        RECT 47.490 118.275 48.330 118.445 ;
        RECT 48.780 118.275 49.620 118.445 ;
        RECT 50.070 118.275 50.910 118.445 ;
        RECT 51.360 118.275 52.200 118.445 ;
        RECT 52.650 118.275 53.490 118.445 ;
        RECT 38.150 117.725 38.320 118.025 ;
        RECT 39.440 117.725 39.610 118.025 ;
        RECT 40.730 117.725 40.900 118.025 ;
        RECT 42.020 117.725 42.190 118.025 ;
        RECT 43.310 117.725 43.480 118.025 ;
        RECT 44.600 117.725 44.770 118.025 ;
        RECT 45.890 117.725 46.060 118.025 ;
        RECT 47.180 117.725 47.350 118.025 ;
        RECT 48.470 117.725 48.640 118.025 ;
        RECT 49.760 117.725 49.930 118.025 ;
        RECT 51.050 117.725 51.220 118.025 ;
        RECT 52.340 117.725 52.510 118.025 ;
        RECT 53.630 117.725 53.800 118.025 ;
        RECT 35.480 116.940 37.480 117.390 ;
        RECT 38.330 116.840 53.580 117.090 ;
        RECT 55.330 114.990 55.530 124.690 ;
        RECT 30.580 114.790 55.530 114.990 ;
        RECT 56.680 113.340 56.880 126.340 ;
        RECT 29.280 113.140 56.880 113.340 ;
        RECT 128.915 127.990 129.755 128.160 ;
        RECT 130.205 127.990 131.045 128.160 ;
        RECT 128.605 126.815 128.775 127.695 ;
        RECT 129.895 126.815 130.065 127.695 ;
        RECT 131.185 126.815 131.355 127.695 ;
        RECT 58.880 122.840 59.480 124.840 ;
        RECT 57.880 114.940 58.380 117.140 ;
        RECT 48.380 111.740 53.980 112.140 ;
        RECT 48.900 110.850 50.885 111.040 ;
        RECT 54.895 110.850 56.880 111.040 ;
        RECT 59.090 110.860 59.280 112.845 ;
        RECT 65.065 124.985 65.235 125.865 ;
        RECT 66.355 124.985 66.525 125.865 ;
        RECT 67.645 124.985 67.815 125.865 ;
        RECT 132.520 126.790 133.020 127.690 ;
        RECT 68.980 125.040 69.480 125.940 ;
        RECT 65.375 124.565 66.215 124.735 ;
        RECT 66.665 124.565 67.505 124.735 ;
        RECT 65.375 121.340 66.215 121.510 ;
        RECT 66.665 121.340 67.505 121.510 ;
        RECT 65.065 120.165 65.235 121.045 ;
        RECT 66.355 120.165 66.525 121.045 ;
        RECT 67.645 120.165 67.815 121.045 ;
        RECT 68.980 120.140 69.480 121.040 ;
        RECT 65.065 117.685 65.235 118.565 ;
        RECT 66.355 117.685 66.525 118.565 ;
        RECT 67.645 117.685 67.815 118.565 ;
        RECT 68.980 117.740 69.480 118.640 ;
        RECT 65.375 117.265 66.215 117.435 ;
        RECT 66.665 117.265 67.505 117.435 ;
        RECT 63.615 114.015 63.785 114.185 ;
        RECT 64.075 114.015 64.245 114.185 ;
        RECT 64.535 114.015 64.705 114.185 ;
        RECT 64.995 114.015 65.165 114.185 ;
        RECT 65.455 114.015 65.625 114.185 ;
        RECT 65.915 114.015 66.085 114.185 ;
        RECT 66.375 114.015 66.545 114.185 ;
        RECT 66.835 114.015 67.005 114.185 ;
        RECT 67.295 114.015 67.465 114.185 ;
        RECT 67.755 114.015 67.925 114.185 ;
        RECT 68.215 114.015 68.385 114.185 ;
        RECT 64.190 112.490 66.630 112.660 ;
        RECT 67.250 112.160 67.490 112.980 ;
        RECT 92.820 125.690 120.420 125.890 ;
        RECT 92.820 112.690 93.020 125.690 ;
        RECT 94.120 124.040 119.070 124.240 ;
        RECT 94.120 114.340 94.320 124.040 ;
        RECT 99.220 122.190 117.120 122.390 ;
        RECT 101.690 120.810 101.860 121.690 ;
        RECT 102.980 120.810 103.150 121.690 ;
        RECT 104.270 120.810 104.440 121.690 ;
        RECT 105.560 120.810 105.730 121.690 ;
        RECT 106.850 120.810 107.020 121.690 ;
        RECT 108.140 120.810 108.310 121.690 ;
        RECT 109.430 120.810 109.600 121.690 ;
        RECT 110.720 120.810 110.890 121.690 ;
        RECT 112.010 120.810 112.180 121.690 ;
        RECT 113.300 120.810 113.470 121.690 ;
        RECT 114.590 120.810 114.760 121.690 ;
        RECT 115.880 120.810 116.050 121.690 ;
        RECT 117.170 120.810 117.340 121.690 ;
        RECT 102.000 120.345 102.840 120.515 ;
        RECT 103.290 120.345 104.130 120.515 ;
        RECT 104.580 120.345 105.420 120.515 ;
        RECT 105.870 120.345 106.710 120.515 ;
        RECT 107.160 120.345 108.000 120.515 ;
        RECT 108.450 120.345 109.290 120.515 ;
        RECT 109.740 120.345 110.580 120.515 ;
        RECT 111.030 120.345 111.870 120.515 ;
        RECT 112.320 120.345 113.160 120.515 ;
        RECT 113.610 120.345 114.450 120.515 ;
        RECT 114.900 120.345 115.740 120.515 ;
        RECT 116.190 120.345 117.030 120.515 ;
        RECT 103.290 119.805 104.130 119.975 ;
        RECT 107.160 119.805 108.000 119.975 ;
        RECT 108.450 119.805 109.290 119.975 ;
        RECT 112.320 119.805 113.160 119.975 ;
        RECT 113.610 119.805 114.450 119.975 ;
        RECT 101.690 118.675 101.860 119.555 ;
        RECT 102.980 118.675 103.150 119.555 ;
        RECT 104.270 118.675 104.440 119.555 ;
        RECT 105.560 118.675 105.730 119.555 ;
        RECT 106.850 118.675 107.020 119.555 ;
        RECT 108.140 118.675 108.310 119.555 ;
        RECT 109.430 118.675 109.600 119.555 ;
        RECT 110.720 118.675 110.890 119.555 ;
        RECT 112.010 118.675 112.180 119.555 ;
        RECT 113.300 118.675 113.470 119.555 ;
        RECT 114.590 118.675 114.760 119.555 ;
        RECT 115.880 118.675 116.050 119.555 ;
        RECT 117.170 118.675 117.340 119.555 ;
        RECT 102.000 118.255 102.840 118.425 ;
        RECT 104.580 118.255 105.420 118.425 ;
        RECT 105.870 118.255 106.710 118.425 ;
        RECT 109.740 118.255 110.580 118.425 ;
        RECT 111.030 118.255 111.870 118.425 ;
        RECT 114.900 118.255 115.740 118.425 ;
        RECT 116.190 118.255 117.030 118.425 ;
        RECT 102.000 117.625 102.840 117.795 ;
        RECT 103.290 117.625 104.130 117.795 ;
        RECT 104.580 117.625 105.420 117.795 ;
        RECT 105.870 117.625 106.710 117.795 ;
        RECT 107.160 117.625 108.000 117.795 ;
        RECT 108.450 117.625 109.290 117.795 ;
        RECT 109.740 117.625 110.580 117.795 ;
        RECT 111.030 117.625 111.870 117.795 ;
        RECT 112.320 117.625 113.160 117.795 ;
        RECT 113.610 117.625 114.450 117.795 ;
        RECT 114.900 117.625 115.740 117.795 ;
        RECT 116.190 117.625 117.030 117.795 ;
        RECT 101.690 117.075 101.860 117.375 ;
        RECT 102.980 117.075 103.150 117.375 ;
        RECT 104.270 117.075 104.440 117.375 ;
        RECT 105.560 117.075 105.730 117.375 ;
        RECT 106.850 117.075 107.020 117.375 ;
        RECT 108.140 117.075 108.310 117.375 ;
        RECT 109.430 117.075 109.600 117.375 ;
        RECT 110.720 117.075 110.890 117.375 ;
        RECT 112.010 117.075 112.180 117.375 ;
        RECT 113.300 117.075 113.470 117.375 ;
        RECT 114.590 117.075 114.760 117.375 ;
        RECT 115.880 117.075 116.050 117.375 ;
        RECT 117.170 117.075 117.340 117.375 ;
        RECT 99.020 116.290 101.020 116.740 ;
        RECT 101.870 116.190 117.120 116.440 ;
        RECT 118.870 114.340 119.070 124.040 ;
        RECT 94.120 114.140 119.070 114.340 ;
        RECT 120.220 112.690 120.420 125.690 ;
        RECT 92.820 112.490 120.420 112.690 ;
        RECT 122.420 122.190 123.020 124.190 ;
        RECT 121.420 114.290 121.920 116.490 ;
        RECT 63.615 111.295 63.785 111.465 ;
        RECT 64.075 111.295 64.245 111.465 ;
        RECT 64.535 111.295 64.705 111.465 ;
        RECT 64.995 111.295 65.165 111.465 ;
        RECT 65.455 111.295 65.625 111.465 ;
        RECT 65.915 111.295 66.085 111.465 ;
        RECT 66.375 111.295 66.545 111.465 ;
        RECT 66.835 111.295 67.005 111.465 ;
        RECT 67.295 111.295 67.465 111.465 ;
        RECT 67.755 111.295 67.925 111.465 ;
        RECT 68.215 111.295 68.385 111.465 ;
        RECT 111.920 111.090 117.520 111.490 ;
        RECT 112.440 110.200 114.425 110.390 ;
        RECT 118.435 110.200 120.420 110.390 ;
        RECT 122.630 110.210 122.820 112.195 ;
        RECT 128.605 124.335 128.775 125.215 ;
        RECT 129.895 124.335 130.065 125.215 ;
        RECT 131.185 124.335 131.355 125.215 ;
        RECT 132.520 124.390 133.020 125.290 ;
        RECT 128.915 123.915 129.755 124.085 ;
        RECT 130.205 123.915 131.045 124.085 ;
        RECT 128.915 120.690 129.755 120.860 ;
        RECT 130.205 120.690 131.045 120.860 ;
        RECT 128.605 119.515 128.775 120.395 ;
        RECT 129.895 119.515 130.065 120.395 ;
        RECT 131.185 119.515 131.355 120.395 ;
        RECT 132.520 119.490 133.020 120.390 ;
        RECT 128.605 117.035 128.775 117.915 ;
        RECT 129.895 117.035 130.065 117.915 ;
        RECT 131.185 117.035 131.355 117.915 ;
        RECT 132.520 117.090 133.020 117.990 ;
        RECT 128.915 116.615 129.755 116.785 ;
        RECT 130.205 116.615 131.045 116.785 ;
        RECT 127.155 113.365 127.325 113.535 ;
        RECT 127.615 113.365 127.785 113.535 ;
        RECT 128.075 113.365 128.245 113.535 ;
        RECT 128.535 113.365 128.705 113.535 ;
        RECT 128.995 113.365 129.165 113.535 ;
        RECT 129.455 113.365 129.625 113.535 ;
        RECT 129.915 113.365 130.085 113.535 ;
        RECT 130.375 113.365 130.545 113.535 ;
        RECT 130.835 113.365 131.005 113.535 ;
        RECT 131.295 113.365 131.465 113.535 ;
        RECT 131.755 113.365 131.925 113.535 ;
        RECT 127.730 111.840 130.170 112.010 ;
        RECT 130.790 111.510 131.030 112.330 ;
        RECT 127.155 110.645 127.325 110.815 ;
        RECT 127.615 110.645 127.785 110.815 ;
        RECT 128.075 110.645 128.245 110.815 ;
        RECT 128.535 110.645 128.705 110.815 ;
        RECT 128.995 110.645 129.165 110.815 ;
        RECT 129.455 110.645 129.625 110.815 ;
        RECT 129.915 110.645 130.085 110.815 ;
        RECT 130.375 110.645 130.545 110.815 ;
        RECT 130.835 110.645 131.005 110.815 ;
        RECT 131.295 110.645 131.465 110.815 ;
        RECT 131.755 110.645 131.925 110.815 ;
        RECT 64.755 93.410 65.595 93.580 ;
        RECT 66.045 93.410 66.885 93.580 ;
        RECT 64.445 92.235 64.615 93.115 ;
        RECT 65.735 92.235 65.905 93.115 ;
        RECT 67.025 92.235 67.195 93.115 ;
        RECT 68.360 92.210 68.860 93.110 ;
        RECT 28.660 91.110 56.260 91.310 ;
        RECT 28.660 78.110 28.860 91.110 ;
        RECT 29.960 89.460 54.910 89.660 ;
        RECT 29.960 79.760 30.160 89.460 ;
        RECT 35.060 87.610 52.960 87.810 ;
        RECT 37.530 86.230 37.700 87.110 ;
        RECT 38.820 86.230 38.990 87.110 ;
        RECT 40.110 86.230 40.280 87.110 ;
        RECT 41.400 86.230 41.570 87.110 ;
        RECT 42.690 86.230 42.860 87.110 ;
        RECT 43.980 86.230 44.150 87.110 ;
        RECT 45.270 86.230 45.440 87.110 ;
        RECT 46.560 86.230 46.730 87.110 ;
        RECT 47.850 86.230 48.020 87.110 ;
        RECT 49.140 86.230 49.310 87.110 ;
        RECT 50.430 86.230 50.600 87.110 ;
        RECT 51.720 86.230 51.890 87.110 ;
        RECT 53.010 86.230 53.180 87.110 ;
        RECT 37.840 85.765 38.680 85.935 ;
        RECT 39.130 85.765 39.970 85.935 ;
        RECT 40.420 85.765 41.260 85.935 ;
        RECT 41.710 85.765 42.550 85.935 ;
        RECT 43.000 85.765 43.840 85.935 ;
        RECT 44.290 85.765 45.130 85.935 ;
        RECT 45.580 85.765 46.420 85.935 ;
        RECT 46.870 85.765 47.710 85.935 ;
        RECT 48.160 85.765 49.000 85.935 ;
        RECT 49.450 85.765 50.290 85.935 ;
        RECT 50.740 85.765 51.580 85.935 ;
        RECT 52.030 85.765 52.870 85.935 ;
        RECT 39.130 85.225 39.970 85.395 ;
        RECT 43.000 85.225 43.840 85.395 ;
        RECT 44.290 85.225 45.130 85.395 ;
        RECT 48.160 85.225 49.000 85.395 ;
        RECT 49.450 85.225 50.290 85.395 ;
        RECT 37.530 84.095 37.700 84.975 ;
        RECT 38.820 84.095 38.990 84.975 ;
        RECT 40.110 84.095 40.280 84.975 ;
        RECT 41.400 84.095 41.570 84.975 ;
        RECT 42.690 84.095 42.860 84.975 ;
        RECT 43.980 84.095 44.150 84.975 ;
        RECT 45.270 84.095 45.440 84.975 ;
        RECT 46.560 84.095 46.730 84.975 ;
        RECT 47.850 84.095 48.020 84.975 ;
        RECT 49.140 84.095 49.310 84.975 ;
        RECT 50.430 84.095 50.600 84.975 ;
        RECT 51.720 84.095 51.890 84.975 ;
        RECT 53.010 84.095 53.180 84.975 ;
        RECT 37.840 83.675 38.680 83.845 ;
        RECT 40.420 83.675 41.260 83.845 ;
        RECT 41.710 83.675 42.550 83.845 ;
        RECT 45.580 83.675 46.420 83.845 ;
        RECT 46.870 83.675 47.710 83.845 ;
        RECT 50.740 83.675 51.580 83.845 ;
        RECT 52.030 83.675 52.870 83.845 ;
        RECT 37.840 83.045 38.680 83.215 ;
        RECT 39.130 83.045 39.970 83.215 ;
        RECT 40.420 83.045 41.260 83.215 ;
        RECT 41.710 83.045 42.550 83.215 ;
        RECT 43.000 83.045 43.840 83.215 ;
        RECT 44.290 83.045 45.130 83.215 ;
        RECT 45.580 83.045 46.420 83.215 ;
        RECT 46.870 83.045 47.710 83.215 ;
        RECT 48.160 83.045 49.000 83.215 ;
        RECT 49.450 83.045 50.290 83.215 ;
        RECT 50.740 83.045 51.580 83.215 ;
        RECT 52.030 83.045 52.870 83.215 ;
        RECT 37.530 82.495 37.700 82.795 ;
        RECT 38.820 82.495 38.990 82.795 ;
        RECT 40.110 82.495 40.280 82.795 ;
        RECT 41.400 82.495 41.570 82.795 ;
        RECT 42.690 82.495 42.860 82.795 ;
        RECT 43.980 82.495 44.150 82.795 ;
        RECT 45.270 82.495 45.440 82.795 ;
        RECT 46.560 82.495 46.730 82.795 ;
        RECT 47.850 82.495 48.020 82.795 ;
        RECT 49.140 82.495 49.310 82.795 ;
        RECT 50.430 82.495 50.600 82.795 ;
        RECT 51.720 82.495 51.890 82.795 ;
        RECT 53.010 82.495 53.180 82.795 ;
        RECT 34.860 81.710 36.860 82.160 ;
        RECT 37.710 81.610 52.960 81.860 ;
        RECT 54.710 79.760 54.910 89.460 ;
        RECT 29.960 79.560 54.910 79.760 ;
        RECT 56.060 78.110 56.260 91.110 ;
        RECT 28.660 77.910 56.260 78.110 ;
        RECT 130.665 92.760 131.505 92.930 ;
        RECT 131.955 92.760 132.795 92.930 ;
        RECT 130.355 91.585 130.525 92.465 ;
        RECT 131.645 91.585 131.815 92.465 ;
        RECT 132.935 91.585 133.105 92.465 ;
        RECT 58.260 87.610 58.860 89.610 ;
        RECT 57.260 79.710 57.760 81.910 ;
        RECT 47.760 76.510 53.360 76.910 ;
        RECT 48.280 75.620 50.265 75.810 ;
        RECT 54.275 75.620 56.260 75.810 ;
        RECT 58.470 75.630 58.660 77.615 ;
        RECT 64.445 89.755 64.615 90.635 ;
        RECT 65.735 89.755 65.905 90.635 ;
        RECT 67.025 89.755 67.195 90.635 ;
        RECT 134.270 91.560 134.770 92.460 ;
        RECT 68.360 89.810 68.860 90.710 ;
        RECT 64.755 89.335 65.595 89.505 ;
        RECT 66.045 89.335 66.885 89.505 ;
        RECT 64.755 86.110 65.595 86.280 ;
        RECT 66.045 86.110 66.885 86.280 ;
        RECT 64.445 84.935 64.615 85.815 ;
        RECT 65.735 84.935 65.905 85.815 ;
        RECT 67.025 84.935 67.195 85.815 ;
        RECT 68.360 84.910 68.860 85.810 ;
        RECT 64.445 82.455 64.615 83.335 ;
        RECT 65.735 82.455 65.905 83.335 ;
        RECT 67.025 82.455 67.195 83.335 ;
        RECT 68.360 82.510 68.860 83.410 ;
        RECT 64.755 82.035 65.595 82.205 ;
        RECT 66.045 82.035 66.885 82.205 ;
        RECT 62.995 78.785 63.165 78.955 ;
        RECT 63.455 78.785 63.625 78.955 ;
        RECT 63.915 78.785 64.085 78.955 ;
        RECT 64.375 78.785 64.545 78.955 ;
        RECT 64.835 78.785 65.005 78.955 ;
        RECT 65.295 78.785 65.465 78.955 ;
        RECT 65.755 78.785 65.925 78.955 ;
        RECT 66.215 78.785 66.385 78.955 ;
        RECT 66.675 78.785 66.845 78.955 ;
        RECT 67.135 78.785 67.305 78.955 ;
        RECT 67.595 78.785 67.765 78.955 ;
        RECT 63.570 77.260 66.010 77.430 ;
        RECT 66.630 76.930 66.870 77.750 ;
        RECT 94.570 90.460 122.170 90.660 ;
        RECT 94.570 77.460 94.770 90.460 ;
        RECT 95.870 88.810 120.820 89.010 ;
        RECT 95.870 79.110 96.070 88.810 ;
        RECT 100.970 86.960 118.870 87.160 ;
        RECT 103.440 85.580 103.610 86.460 ;
        RECT 104.730 85.580 104.900 86.460 ;
        RECT 106.020 85.580 106.190 86.460 ;
        RECT 107.310 85.580 107.480 86.460 ;
        RECT 108.600 85.580 108.770 86.460 ;
        RECT 109.890 85.580 110.060 86.460 ;
        RECT 111.180 85.580 111.350 86.460 ;
        RECT 112.470 85.580 112.640 86.460 ;
        RECT 113.760 85.580 113.930 86.460 ;
        RECT 115.050 85.580 115.220 86.460 ;
        RECT 116.340 85.580 116.510 86.460 ;
        RECT 117.630 85.580 117.800 86.460 ;
        RECT 118.920 85.580 119.090 86.460 ;
        RECT 103.750 85.115 104.590 85.285 ;
        RECT 105.040 85.115 105.880 85.285 ;
        RECT 106.330 85.115 107.170 85.285 ;
        RECT 107.620 85.115 108.460 85.285 ;
        RECT 108.910 85.115 109.750 85.285 ;
        RECT 110.200 85.115 111.040 85.285 ;
        RECT 111.490 85.115 112.330 85.285 ;
        RECT 112.780 85.115 113.620 85.285 ;
        RECT 114.070 85.115 114.910 85.285 ;
        RECT 115.360 85.115 116.200 85.285 ;
        RECT 116.650 85.115 117.490 85.285 ;
        RECT 117.940 85.115 118.780 85.285 ;
        RECT 105.040 84.575 105.880 84.745 ;
        RECT 108.910 84.575 109.750 84.745 ;
        RECT 110.200 84.575 111.040 84.745 ;
        RECT 114.070 84.575 114.910 84.745 ;
        RECT 115.360 84.575 116.200 84.745 ;
        RECT 103.440 83.445 103.610 84.325 ;
        RECT 104.730 83.445 104.900 84.325 ;
        RECT 106.020 83.445 106.190 84.325 ;
        RECT 107.310 83.445 107.480 84.325 ;
        RECT 108.600 83.445 108.770 84.325 ;
        RECT 109.890 83.445 110.060 84.325 ;
        RECT 111.180 83.445 111.350 84.325 ;
        RECT 112.470 83.445 112.640 84.325 ;
        RECT 113.760 83.445 113.930 84.325 ;
        RECT 115.050 83.445 115.220 84.325 ;
        RECT 116.340 83.445 116.510 84.325 ;
        RECT 117.630 83.445 117.800 84.325 ;
        RECT 118.920 83.445 119.090 84.325 ;
        RECT 103.750 83.025 104.590 83.195 ;
        RECT 106.330 83.025 107.170 83.195 ;
        RECT 107.620 83.025 108.460 83.195 ;
        RECT 111.490 83.025 112.330 83.195 ;
        RECT 112.780 83.025 113.620 83.195 ;
        RECT 116.650 83.025 117.490 83.195 ;
        RECT 117.940 83.025 118.780 83.195 ;
        RECT 103.750 82.395 104.590 82.565 ;
        RECT 105.040 82.395 105.880 82.565 ;
        RECT 106.330 82.395 107.170 82.565 ;
        RECT 107.620 82.395 108.460 82.565 ;
        RECT 108.910 82.395 109.750 82.565 ;
        RECT 110.200 82.395 111.040 82.565 ;
        RECT 111.490 82.395 112.330 82.565 ;
        RECT 112.780 82.395 113.620 82.565 ;
        RECT 114.070 82.395 114.910 82.565 ;
        RECT 115.360 82.395 116.200 82.565 ;
        RECT 116.650 82.395 117.490 82.565 ;
        RECT 117.940 82.395 118.780 82.565 ;
        RECT 103.440 81.845 103.610 82.145 ;
        RECT 104.730 81.845 104.900 82.145 ;
        RECT 106.020 81.845 106.190 82.145 ;
        RECT 107.310 81.845 107.480 82.145 ;
        RECT 108.600 81.845 108.770 82.145 ;
        RECT 109.890 81.845 110.060 82.145 ;
        RECT 111.180 81.845 111.350 82.145 ;
        RECT 112.470 81.845 112.640 82.145 ;
        RECT 113.760 81.845 113.930 82.145 ;
        RECT 115.050 81.845 115.220 82.145 ;
        RECT 116.340 81.845 116.510 82.145 ;
        RECT 117.630 81.845 117.800 82.145 ;
        RECT 118.920 81.845 119.090 82.145 ;
        RECT 100.770 81.060 102.770 81.510 ;
        RECT 103.620 80.960 118.870 81.210 ;
        RECT 120.620 79.110 120.820 88.810 ;
        RECT 95.870 78.910 120.820 79.110 ;
        RECT 121.970 77.460 122.170 90.460 ;
        RECT 94.570 77.260 122.170 77.460 ;
        RECT 124.170 86.960 124.770 88.960 ;
        RECT 123.170 79.060 123.670 81.260 ;
        RECT 62.995 76.065 63.165 76.235 ;
        RECT 63.455 76.065 63.625 76.235 ;
        RECT 63.915 76.065 64.085 76.235 ;
        RECT 64.375 76.065 64.545 76.235 ;
        RECT 64.835 76.065 65.005 76.235 ;
        RECT 65.295 76.065 65.465 76.235 ;
        RECT 65.755 76.065 65.925 76.235 ;
        RECT 66.215 76.065 66.385 76.235 ;
        RECT 66.675 76.065 66.845 76.235 ;
        RECT 67.135 76.065 67.305 76.235 ;
        RECT 67.595 76.065 67.765 76.235 ;
        RECT 113.670 75.860 119.270 76.260 ;
        RECT 114.190 74.970 116.175 75.160 ;
        RECT 120.185 74.970 122.170 75.160 ;
        RECT 124.380 74.980 124.570 76.965 ;
        RECT 130.355 89.105 130.525 89.985 ;
        RECT 131.645 89.105 131.815 89.985 ;
        RECT 132.935 89.105 133.105 89.985 ;
        RECT 134.270 89.160 134.770 90.060 ;
        RECT 130.665 88.685 131.505 88.855 ;
        RECT 131.955 88.685 132.795 88.855 ;
        RECT 130.665 85.460 131.505 85.630 ;
        RECT 131.955 85.460 132.795 85.630 ;
        RECT 130.355 84.285 130.525 85.165 ;
        RECT 131.645 84.285 131.815 85.165 ;
        RECT 132.935 84.285 133.105 85.165 ;
        RECT 134.270 84.260 134.770 85.160 ;
        RECT 130.355 81.805 130.525 82.685 ;
        RECT 131.645 81.805 131.815 82.685 ;
        RECT 132.935 81.805 133.105 82.685 ;
        RECT 134.270 81.860 134.770 82.760 ;
        RECT 130.665 81.385 131.505 81.555 ;
        RECT 131.955 81.385 132.795 81.555 ;
        RECT 128.905 78.135 129.075 78.305 ;
        RECT 129.365 78.135 129.535 78.305 ;
        RECT 129.825 78.135 129.995 78.305 ;
        RECT 130.285 78.135 130.455 78.305 ;
        RECT 130.745 78.135 130.915 78.305 ;
        RECT 131.205 78.135 131.375 78.305 ;
        RECT 131.665 78.135 131.835 78.305 ;
        RECT 132.125 78.135 132.295 78.305 ;
        RECT 132.585 78.135 132.755 78.305 ;
        RECT 133.045 78.135 133.215 78.305 ;
        RECT 133.505 78.135 133.675 78.305 ;
        RECT 129.480 76.610 131.920 76.780 ;
        RECT 132.540 76.280 132.780 77.100 ;
        RECT 128.905 75.415 129.075 75.585 ;
        RECT 129.365 75.415 129.535 75.585 ;
        RECT 129.825 75.415 129.995 75.585 ;
        RECT 130.285 75.415 130.455 75.585 ;
        RECT 130.745 75.415 130.915 75.585 ;
        RECT 131.205 75.415 131.375 75.585 ;
        RECT 131.665 75.415 131.835 75.585 ;
        RECT 132.125 75.415 132.295 75.585 ;
        RECT 132.585 75.415 132.755 75.585 ;
        RECT 133.045 75.415 133.215 75.585 ;
        RECT 133.505 75.415 133.675 75.585 ;
      LAYER met1 ;
        RECT 64.450 191.600 66.750 193.100 ;
        RECT 128.520 192.380 130.820 193.880 ;
        RECT 128.555 192.350 129.515 192.380 ;
        RECT 129.845 192.350 130.805 192.380 ;
        RECT 133.120 192.180 137.320 192.380 ;
        RECT 64.485 191.570 65.445 191.600 ;
        RECT 65.775 191.570 66.735 191.600 ;
        RECT 69.050 191.400 73.250 191.600 ;
        RECT 63.350 190.300 64.650 191.400 ;
        RECT 65.350 189.900 65.850 191.400 ;
        RECT 66.550 190.300 67.850 191.400 ;
        RECT 68.050 190.300 73.250 191.400 ;
        RECT 127.420 191.080 128.720 192.180 ;
        RECT 129.420 190.680 129.920 192.180 ;
        RECT 130.620 191.080 131.920 192.180 ;
        RECT 132.120 191.080 137.320 192.180 ;
        RECT 133.120 190.880 137.320 191.080 ;
        RECT 69.050 190.100 73.250 190.300 ;
        RECT 27.950 188.800 56.450 189.800 ;
        RECT 64.050 189.500 67.150 189.900 ;
        RECT 64.050 189.000 64.550 189.500 ;
        RECT 66.650 189.000 67.150 189.500 ;
        RECT 92.020 189.580 120.520 190.580 ;
        RECT 128.120 190.280 131.220 190.680 ;
        RECT 128.120 189.780 128.620 190.280 ;
        RECT 130.720 189.780 131.220 190.280 ;
        RECT 133.120 189.780 137.320 189.980 ;
        RECT 69.050 189.000 73.250 189.200 ;
        RECT 27.950 176.800 28.950 188.800 ;
        RECT 29.450 187.300 54.950 188.300 ;
        RECT 29.450 178.300 30.450 187.300 ;
        RECT 34.550 185.600 53.000 186.200 ;
        RECT 37.300 185.360 37.600 185.600 ;
        RECT 37.290 184.360 37.600 185.360 ;
        RECT 38.550 185.350 38.850 185.400 ;
        RECT 38.350 184.400 39.100 185.350 ;
        RECT 39.650 184.400 40.300 185.600 ;
        RECT 41.160 185.350 41.390 185.360 ;
        RECT 40.950 184.400 41.600 185.350 ;
        RECT 42.250 184.400 42.900 185.600 ;
        RECT 37.300 184.155 37.600 184.360 ;
        RECT 38.550 184.350 39.100 184.400 ;
        RECT 39.870 184.360 40.100 184.400 ;
        RECT 41.160 184.360 41.390 184.400 ;
        RECT 42.450 184.360 42.680 184.400 ;
        RECT 38.850 184.155 39.100 184.350 ;
        RECT 43.500 184.155 44.150 185.400 ;
        RECT 44.800 184.400 45.450 185.600 ;
        RECT 46.320 185.350 46.550 185.360 ;
        RECT 46.100 184.400 46.750 185.350 ;
        RECT 47.400 184.400 48.050 185.600 ;
        RECT 45.030 184.360 45.260 184.400 ;
        RECT 46.320 184.360 46.550 184.400 ;
        RECT 47.610 184.360 47.840 184.400 ;
        RECT 48.700 184.155 49.350 185.400 ;
        RECT 50.000 184.400 50.650 185.600 ;
        RECT 52.800 185.360 53.000 185.600 ;
        RECT 51.480 185.350 51.710 185.360 ;
        RECT 51.250 184.400 51.900 185.350 ;
        RECT 50.190 184.360 50.420 184.400 ;
        RECT 51.480 184.360 51.710 184.400 ;
        RECT 52.770 184.360 53.000 185.360 ;
        RECT 52.800 184.200 53.000 184.360 ;
        RECT 37.300 184.150 38.530 184.155 ;
        RECT 37.300 183.950 38.550 184.150 ;
        RECT 38.850 184.125 39.820 184.155 ;
        RECT 40.150 184.125 41.110 184.155 ;
        RECT 41.440 184.125 42.400 184.155 ;
        RECT 42.730 184.125 44.980 184.155 ;
        RECT 45.310 184.125 46.270 184.155 ;
        RECT 46.600 184.125 47.560 184.155 ;
        RECT 47.890 184.125 50.140 184.155 ;
        RECT 50.470 184.125 51.430 184.155 ;
        RECT 38.840 183.955 51.450 184.125 ;
        RECT 38.850 183.950 39.820 183.955 ;
        RECT 37.570 183.925 38.530 183.950 ;
        RECT 38.860 183.925 39.820 183.950 ;
        RECT 40.150 183.925 41.110 183.955 ;
        RECT 41.440 183.925 42.400 183.955 ;
        RECT 42.730 183.925 43.690 183.955 ;
        RECT 44.020 183.925 44.980 183.955 ;
        RECT 45.310 183.925 46.270 183.955 ;
        RECT 46.600 183.925 47.560 183.955 ;
        RECT 47.890 183.925 48.850 183.955 ;
        RECT 49.180 183.925 50.140 183.955 ;
        RECT 50.470 183.925 51.430 183.955 ;
        RECT 51.750 183.950 53.000 184.200 ;
        RECT 51.760 183.925 52.720 183.950 ;
        RECT 38.860 183.585 39.820 183.615 ;
        RECT 40.250 183.585 40.800 183.750 ;
        RECT 42.730 183.585 43.690 183.615 ;
        RECT 44.020 183.585 44.980 183.615 ;
        RECT 47.890 183.585 48.850 183.615 ;
        RECT 49.180 183.585 50.140 183.615 ;
        RECT 38.840 183.415 50.160 183.585 ;
        RECT 38.860 183.385 39.820 183.415 ;
        RECT 37.300 183.225 37.550 183.250 ;
        RECT 37.290 182.225 37.550 183.225 ;
        RECT 38.580 183.200 38.810 183.225 ;
        RECT 38.350 182.250 39.000 183.200 ;
        RECT 39.870 182.700 40.100 183.225 ;
        RECT 40.250 182.850 40.800 183.415 ;
        RECT 42.730 183.385 43.690 183.415 ;
        RECT 44.020 183.385 44.980 183.415 ;
        RECT 47.890 183.385 48.850 183.415 ;
        RECT 49.180 183.385 50.140 183.415 ;
        RECT 41.160 183.200 41.390 183.225 ;
        RECT 42.450 183.200 42.680 183.225 ;
        RECT 43.740 183.200 43.970 183.225 ;
        RECT 45.030 183.200 45.260 183.225 ;
        RECT 46.320 183.200 46.550 183.225 ;
        RECT 47.610 183.200 47.840 183.225 ;
        RECT 48.900 183.200 49.130 183.225 ;
        RECT 39.650 182.250 40.300 182.700 ;
        RECT 40.950 182.250 41.600 183.200 ;
        RECT 42.250 182.250 42.900 183.200 ;
        RECT 43.500 182.250 44.150 183.200 ;
        RECT 44.850 182.250 45.500 183.200 ;
        RECT 46.100 182.250 46.750 183.200 ;
        RECT 47.400 182.250 48.050 183.200 ;
        RECT 48.700 182.250 49.350 183.200 ;
        RECT 50.190 182.650 50.420 183.225 ;
        RECT 50.600 182.800 51.100 183.750 ;
        RECT 51.480 183.200 51.710 183.225 ;
        RECT 49.950 182.250 50.600 182.650 ;
        RECT 38.580 182.225 38.810 182.250 ;
        RECT 39.870 182.225 40.100 182.250 ;
        RECT 41.160 182.225 41.390 182.250 ;
        RECT 42.450 182.225 42.680 182.250 ;
        RECT 43.740 182.225 43.970 182.250 ;
        RECT 45.030 182.225 45.260 182.250 ;
        RECT 46.320 182.225 46.550 182.250 ;
        RECT 47.610 182.225 47.840 182.250 ;
        RECT 48.900 182.225 49.130 182.250 ;
        RECT 50.190 182.225 50.420 182.250 ;
        RECT 37.300 182.200 37.550 182.225 ;
        RECT 37.300 182.065 37.650 182.200 ;
        RECT 50.750 182.065 51.100 182.800 ;
        RECT 51.250 182.250 51.900 183.200 ;
        RECT 51.480 182.225 51.710 182.250 ;
        RECT 52.750 182.200 53.000 183.250 ;
        RECT 52.600 182.065 53.000 182.200 ;
        RECT 37.300 182.050 38.530 182.065 ;
        RECT 37.300 181.550 38.550 182.050 ;
        RECT 40.150 182.035 41.110 182.065 ;
        RECT 41.440 182.035 42.400 182.065 ;
        RECT 45.310 182.035 46.270 182.065 ;
        RECT 46.600 182.035 47.560 182.065 ;
        RECT 50.470 182.035 51.430 182.065 ;
        RECT 51.760 182.050 53.000 182.065 ;
        RECT 40.130 181.865 51.450 182.035 ;
        RECT 40.150 181.835 41.110 181.865 ;
        RECT 41.440 181.835 42.400 181.865 ;
        RECT 45.310 181.835 46.270 181.865 ;
        RECT 46.600 181.835 47.560 181.865 ;
        RECT 50.470 181.835 51.430 181.865 ;
        RECT 37.300 181.150 41.150 181.550 ;
        RECT 44.550 181.500 45.750 181.650 ;
        RECT 51.700 181.550 53.000 182.050 ;
        RECT 41.400 181.200 48.900 181.500 ;
        RECT 44.550 181.150 45.750 181.200 ;
        RECT 37.300 181.050 41.250 181.150 ;
        RECT 37.300 181.045 41.370 181.050 ;
        RECT 37.290 180.625 41.390 181.045 ;
        RECT 42.350 180.625 42.800 181.050 ;
        RECT 34.550 179.800 36.750 180.500 ;
        RECT 37.300 180.200 41.370 180.625 ;
        RECT 43.500 180.200 44.200 181.050 ;
        RECT 44.925 180.600 45.375 181.150 ;
        RECT 49.150 181.050 53.000 181.550 ;
        RECT 46.100 180.200 46.800 181.050 ;
        RECT 47.525 180.625 47.900 181.050 ;
        RECT 48.900 180.200 53.000 181.050 ;
        RECT 37.300 179.650 53.000 180.200 ;
        RECT 53.950 178.300 54.950 187.300 ;
        RECT 29.450 177.300 54.950 178.300 ;
        RECT 55.450 176.800 56.450 188.800 ;
        RECT 57.750 185.600 59.050 188.200 ;
        RECT 63.350 187.900 64.650 189.000 ;
        RECT 64.205 187.885 64.435 187.900 ;
        RECT 65.495 187.885 65.725 188.885 ;
        RECT 66.550 187.900 67.850 189.000 ;
        RECT 68.050 187.900 73.250 189.000 ;
        RECT 66.785 187.885 67.015 187.900 ;
        RECT 64.485 187.700 65.445 187.725 ;
        RECT 65.775 187.700 66.735 187.725 ;
        RECT 69.050 187.700 73.250 187.900 ;
        RECT 64.450 186.200 66.750 187.700 ;
        RECT 64.450 184.300 66.750 185.800 ;
        RECT 64.485 184.270 65.445 184.300 ;
        RECT 65.775 184.270 66.735 184.300 ;
        RECT 69.050 184.100 73.250 184.300 ;
        RECT 63.350 183.000 64.650 184.100 ;
        RECT 65.350 182.600 65.850 184.100 ;
        RECT 66.550 183.000 67.850 184.100 ;
        RECT 68.050 183.000 73.250 184.100 ;
        RECT 69.050 182.800 73.250 183.000 ;
        RECT 64.050 182.200 67.150 182.600 ;
        RECT 64.050 181.700 64.550 182.200 ;
        RECT 66.650 181.700 67.150 182.200 ;
        RECT 69.050 181.700 73.250 181.900 ;
        RECT 63.350 180.600 64.650 181.700 ;
        RECT 64.205 180.585 64.435 180.600 ;
        RECT 65.495 180.585 65.725 181.585 ;
        RECT 66.550 180.600 67.850 181.700 ;
        RECT 68.050 180.600 73.250 181.700 ;
        RECT 66.785 180.585 67.015 180.600 ;
        RECT 64.485 180.400 65.445 180.425 ;
        RECT 65.775 180.400 66.735 180.425 ;
        RECT 69.050 180.400 73.250 180.600 ;
        RECT 56.950 177.800 57.650 180.200 ;
        RECT 64.450 178.900 66.750 180.400 ;
        RECT 92.020 177.580 93.020 189.580 ;
        RECT 93.520 188.080 119.020 189.080 ;
        RECT 93.520 179.080 94.520 188.080 ;
        RECT 98.620 186.380 117.070 186.980 ;
        RECT 101.370 186.140 101.670 186.380 ;
        RECT 101.360 185.140 101.670 186.140 ;
        RECT 102.620 186.130 102.920 186.180 ;
        RECT 102.420 185.180 103.170 186.130 ;
        RECT 103.720 185.180 104.370 186.380 ;
        RECT 105.230 186.130 105.460 186.140 ;
        RECT 105.020 185.180 105.670 186.130 ;
        RECT 106.320 185.180 106.970 186.380 ;
        RECT 101.370 184.935 101.670 185.140 ;
        RECT 102.620 185.130 103.170 185.180 ;
        RECT 103.940 185.140 104.170 185.180 ;
        RECT 105.230 185.140 105.460 185.180 ;
        RECT 106.520 185.140 106.750 185.180 ;
        RECT 102.920 184.935 103.170 185.130 ;
        RECT 107.570 184.935 108.220 186.180 ;
        RECT 108.870 185.180 109.520 186.380 ;
        RECT 110.390 186.130 110.620 186.140 ;
        RECT 110.170 185.180 110.820 186.130 ;
        RECT 111.470 185.180 112.120 186.380 ;
        RECT 109.100 185.140 109.330 185.180 ;
        RECT 110.390 185.140 110.620 185.180 ;
        RECT 111.680 185.140 111.910 185.180 ;
        RECT 112.770 184.935 113.420 186.180 ;
        RECT 114.070 185.180 114.720 186.380 ;
        RECT 116.870 186.140 117.070 186.380 ;
        RECT 115.550 186.130 115.780 186.140 ;
        RECT 115.320 185.180 115.970 186.130 ;
        RECT 114.260 185.140 114.490 185.180 ;
        RECT 115.550 185.140 115.780 185.180 ;
        RECT 116.840 185.140 117.070 186.140 ;
        RECT 116.870 184.980 117.070 185.140 ;
        RECT 101.370 184.930 102.600 184.935 ;
        RECT 101.370 184.730 102.620 184.930 ;
        RECT 102.920 184.905 103.890 184.935 ;
        RECT 104.220 184.905 105.180 184.935 ;
        RECT 105.510 184.905 106.470 184.935 ;
        RECT 106.800 184.905 109.050 184.935 ;
        RECT 109.380 184.905 110.340 184.935 ;
        RECT 110.670 184.905 111.630 184.935 ;
        RECT 111.960 184.905 114.210 184.935 ;
        RECT 114.540 184.905 115.500 184.935 ;
        RECT 102.910 184.735 115.520 184.905 ;
        RECT 102.920 184.730 103.890 184.735 ;
        RECT 101.640 184.705 102.600 184.730 ;
        RECT 102.930 184.705 103.890 184.730 ;
        RECT 104.220 184.705 105.180 184.735 ;
        RECT 105.510 184.705 106.470 184.735 ;
        RECT 106.800 184.705 107.760 184.735 ;
        RECT 108.090 184.705 109.050 184.735 ;
        RECT 109.380 184.705 110.340 184.735 ;
        RECT 110.670 184.705 111.630 184.735 ;
        RECT 111.960 184.705 112.920 184.735 ;
        RECT 113.250 184.705 114.210 184.735 ;
        RECT 114.540 184.705 115.500 184.735 ;
        RECT 115.820 184.730 117.070 184.980 ;
        RECT 115.830 184.705 116.790 184.730 ;
        RECT 102.930 184.365 103.890 184.395 ;
        RECT 104.320 184.365 104.870 184.530 ;
        RECT 106.800 184.365 107.760 184.395 ;
        RECT 108.090 184.365 109.050 184.395 ;
        RECT 111.960 184.365 112.920 184.395 ;
        RECT 113.250 184.365 114.210 184.395 ;
        RECT 102.910 184.195 114.230 184.365 ;
        RECT 102.930 184.165 103.890 184.195 ;
        RECT 101.370 184.005 101.620 184.030 ;
        RECT 101.360 183.005 101.620 184.005 ;
        RECT 102.650 183.980 102.880 184.005 ;
        RECT 102.420 183.030 103.070 183.980 ;
        RECT 103.940 183.480 104.170 184.005 ;
        RECT 104.320 183.630 104.870 184.195 ;
        RECT 106.800 184.165 107.760 184.195 ;
        RECT 108.090 184.165 109.050 184.195 ;
        RECT 111.960 184.165 112.920 184.195 ;
        RECT 113.250 184.165 114.210 184.195 ;
        RECT 105.230 183.980 105.460 184.005 ;
        RECT 106.520 183.980 106.750 184.005 ;
        RECT 107.810 183.980 108.040 184.005 ;
        RECT 109.100 183.980 109.330 184.005 ;
        RECT 110.390 183.980 110.620 184.005 ;
        RECT 111.680 183.980 111.910 184.005 ;
        RECT 112.970 183.980 113.200 184.005 ;
        RECT 103.720 183.030 104.370 183.480 ;
        RECT 105.020 183.030 105.670 183.980 ;
        RECT 106.320 183.030 106.970 183.980 ;
        RECT 107.570 183.030 108.220 183.980 ;
        RECT 108.920 183.030 109.570 183.980 ;
        RECT 110.170 183.030 110.820 183.980 ;
        RECT 111.470 183.030 112.120 183.980 ;
        RECT 112.770 183.030 113.420 183.980 ;
        RECT 114.260 183.430 114.490 184.005 ;
        RECT 114.670 183.580 115.170 184.530 ;
        RECT 115.550 183.980 115.780 184.005 ;
        RECT 114.020 183.030 114.670 183.430 ;
        RECT 102.650 183.005 102.880 183.030 ;
        RECT 103.940 183.005 104.170 183.030 ;
        RECT 105.230 183.005 105.460 183.030 ;
        RECT 106.520 183.005 106.750 183.030 ;
        RECT 107.810 183.005 108.040 183.030 ;
        RECT 109.100 183.005 109.330 183.030 ;
        RECT 110.390 183.005 110.620 183.030 ;
        RECT 111.680 183.005 111.910 183.030 ;
        RECT 112.970 183.005 113.200 183.030 ;
        RECT 114.260 183.005 114.490 183.030 ;
        RECT 101.370 182.980 101.620 183.005 ;
        RECT 101.370 182.845 101.720 182.980 ;
        RECT 114.820 182.845 115.170 183.580 ;
        RECT 115.320 183.030 115.970 183.980 ;
        RECT 115.550 183.005 115.780 183.030 ;
        RECT 116.820 182.980 117.070 184.030 ;
        RECT 116.670 182.845 117.070 182.980 ;
        RECT 101.370 182.830 102.600 182.845 ;
        RECT 101.370 182.330 102.620 182.830 ;
        RECT 104.220 182.815 105.180 182.845 ;
        RECT 105.510 182.815 106.470 182.845 ;
        RECT 109.380 182.815 110.340 182.845 ;
        RECT 110.670 182.815 111.630 182.845 ;
        RECT 114.540 182.815 115.500 182.845 ;
        RECT 115.830 182.830 117.070 182.845 ;
        RECT 104.200 182.645 115.520 182.815 ;
        RECT 104.220 182.615 105.180 182.645 ;
        RECT 105.510 182.615 106.470 182.645 ;
        RECT 109.380 182.615 110.340 182.645 ;
        RECT 110.670 182.615 111.630 182.645 ;
        RECT 114.540 182.615 115.500 182.645 ;
        RECT 101.370 181.930 105.220 182.330 ;
        RECT 108.620 182.280 109.820 182.430 ;
        RECT 115.770 182.330 117.070 182.830 ;
        RECT 105.470 181.980 112.970 182.280 ;
        RECT 108.620 181.930 109.820 181.980 ;
        RECT 101.370 181.830 105.320 181.930 ;
        RECT 101.370 181.825 105.440 181.830 ;
        RECT 101.360 181.405 105.460 181.825 ;
        RECT 106.420 181.405 106.870 181.830 ;
        RECT 98.620 180.580 100.820 181.280 ;
        RECT 101.370 180.980 105.440 181.405 ;
        RECT 107.570 180.980 108.270 181.830 ;
        RECT 108.995 181.380 109.445 181.930 ;
        RECT 113.220 181.830 117.070 182.330 ;
        RECT 110.170 180.980 110.870 181.830 ;
        RECT 111.595 181.405 111.970 181.830 ;
        RECT 112.970 180.980 117.070 181.830 ;
        RECT 101.370 180.430 117.070 180.980 ;
        RECT 118.020 179.080 119.020 188.080 ;
        RECT 93.520 178.080 119.020 179.080 ;
        RECT 119.520 177.580 120.520 189.580 ;
        RECT 121.820 186.380 123.120 188.980 ;
        RECT 127.420 188.680 128.720 189.780 ;
        RECT 128.275 188.665 128.505 188.680 ;
        RECT 129.565 188.665 129.795 189.665 ;
        RECT 130.620 188.680 131.920 189.780 ;
        RECT 132.120 188.680 137.320 189.780 ;
        RECT 130.855 188.665 131.085 188.680 ;
        RECT 128.555 188.480 129.515 188.505 ;
        RECT 129.845 188.480 130.805 188.505 ;
        RECT 133.120 188.480 137.320 188.680 ;
        RECT 128.520 186.980 130.820 188.480 ;
        RECT 128.520 185.080 130.820 186.580 ;
        RECT 128.555 185.050 129.515 185.080 ;
        RECT 129.845 185.050 130.805 185.080 ;
        RECT 133.120 184.880 137.320 185.080 ;
        RECT 127.420 183.780 128.720 184.880 ;
        RECT 129.420 183.380 129.920 184.880 ;
        RECT 130.620 183.780 131.920 184.880 ;
        RECT 132.120 183.780 137.320 184.880 ;
        RECT 133.120 183.580 137.320 183.780 ;
        RECT 128.120 182.980 131.220 183.380 ;
        RECT 128.120 182.480 128.620 182.980 ;
        RECT 130.720 182.480 131.220 182.980 ;
        RECT 133.120 182.480 137.320 182.680 ;
        RECT 127.420 181.380 128.720 182.480 ;
        RECT 128.275 181.365 128.505 181.380 ;
        RECT 129.565 181.365 129.795 182.365 ;
        RECT 130.620 181.380 131.920 182.480 ;
        RECT 132.120 181.380 137.320 182.480 ;
        RECT 130.855 181.365 131.085 181.380 ;
        RECT 128.555 181.180 129.515 181.205 ;
        RECT 129.845 181.180 130.805 181.205 ;
        RECT 133.120 181.180 137.320 181.380 ;
        RECT 121.020 178.580 121.720 180.980 ;
        RECT 128.520 179.680 130.820 181.180 ;
        RECT 126.710 177.600 131.770 178.080 ;
        RECT 62.640 176.820 67.700 177.300 ;
        RECT 27.950 175.800 56.450 176.800 ;
        RECT 92.020 176.580 120.520 177.580 ;
        RECT 47.450 174.600 53.250 175.200 ;
        RECT 57.850 174.500 58.850 175.900 ;
        RECT 60.850 175.000 65.850 176.100 ;
        RECT 66.350 175.000 68.350 176.100 ;
        RECT 111.520 175.380 117.320 175.980 ;
        RECT 121.920 175.280 122.920 176.680 ;
        RECT 124.920 175.780 129.920 176.880 ;
        RECT 130.420 175.780 132.420 176.880 ;
        RECT 48.010 173.780 50.115 174.030 ;
        RECT 53.950 173.400 58.850 174.500 ;
        RECT 62.640 174.100 67.700 174.580 ;
        RECT 112.080 174.560 114.185 174.810 ;
        RECT 118.020 174.180 122.920 175.280 ;
        RECT 126.710 174.880 131.770 175.360 ;
        RECT 64.680 162.160 66.980 163.660 ;
        RECT 64.715 162.130 65.675 162.160 ;
        RECT 66.005 162.130 66.965 162.160 ;
        RECT 69.280 161.960 73.480 162.160 ;
        RECT 63.580 160.860 64.880 161.960 ;
        RECT 65.580 160.460 66.080 161.960 ;
        RECT 66.780 160.860 68.080 161.960 ;
        RECT 68.280 160.860 73.480 161.960 ;
        RECT 128.340 161.780 130.640 163.280 ;
        RECT 128.375 161.750 129.335 161.780 ;
        RECT 129.665 161.750 130.625 161.780 ;
        RECT 132.940 161.580 137.140 161.780 ;
        RECT 69.280 160.660 73.480 160.860 ;
        RECT 127.240 160.480 128.540 161.580 ;
        RECT 28.180 159.360 56.680 160.360 ;
        RECT 64.280 160.060 67.380 160.460 ;
        RECT 129.240 160.080 129.740 161.580 ;
        RECT 130.440 160.480 131.740 161.580 ;
        RECT 131.940 160.480 137.140 161.580 ;
        RECT 132.940 160.280 137.140 160.480 ;
        RECT 64.280 159.560 64.780 160.060 ;
        RECT 66.880 159.560 67.380 160.060 ;
        RECT 69.280 159.560 73.480 159.760 ;
        RECT 28.180 147.360 29.180 159.360 ;
        RECT 29.680 157.860 55.180 158.860 ;
        RECT 29.680 148.860 30.680 157.860 ;
        RECT 34.780 156.160 53.230 156.760 ;
        RECT 37.530 155.920 37.830 156.160 ;
        RECT 37.520 154.920 37.830 155.920 ;
        RECT 38.780 155.910 39.080 155.960 ;
        RECT 38.580 154.960 39.330 155.910 ;
        RECT 39.880 154.960 40.530 156.160 ;
        RECT 41.390 155.910 41.620 155.920 ;
        RECT 41.180 154.960 41.830 155.910 ;
        RECT 42.480 154.960 43.130 156.160 ;
        RECT 37.530 154.715 37.830 154.920 ;
        RECT 38.780 154.910 39.330 154.960 ;
        RECT 40.100 154.920 40.330 154.960 ;
        RECT 41.390 154.920 41.620 154.960 ;
        RECT 42.680 154.920 42.910 154.960 ;
        RECT 39.080 154.715 39.330 154.910 ;
        RECT 43.730 154.715 44.380 155.960 ;
        RECT 45.030 154.960 45.680 156.160 ;
        RECT 46.550 155.910 46.780 155.920 ;
        RECT 46.330 154.960 46.980 155.910 ;
        RECT 47.630 154.960 48.280 156.160 ;
        RECT 45.260 154.920 45.490 154.960 ;
        RECT 46.550 154.920 46.780 154.960 ;
        RECT 47.840 154.920 48.070 154.960 ;
        RECT 48.930 154.715 49.580 155.960 ;
        RECT 50.230 154.960 50.880 156.160 ;
        RECT 53.030 155.920 53.230 156.160 ;
        RECT 51.710 155.910 51.940 155.920 ;
        RECT 51.480 154.960 52.130 155.910 ;
        RECT 50.420 154.920 50.650 154.960 ;
        RECT 51.710 154.920 51.940 154.960 ;
        RECT 53.000 154.920 53.230 155.920 ;
        RECT 53.030 154.760 53.230 154.920 ;
        RECT 37.530 154.710 38.760 154.715 ;
        RECT 37.530 154.510 38.780 154.710 ;
        RECT 39.080 154.685 40.050 154.715 ;
        RECT 40.380 154.685 41.340 154.715 ;
        RECT 41.670 154.685 42.630 154.715 ;
        RECT 42.960 154.685 45.210 154.715 ;
        RECT 45.540 154.685 46.500 154.715 ;
        RECT 46.830 154.685 47.790 154.715 ;
        RECT 48.120 154.685 50.370 154.715 ;
        RECT 50.700 154.685 51.660 154.715 ;
        RECT 39.070 154.515 51.680 154.685 ;
        RECT 39.080 154.510 40.050 154.515 ;
        RECT 37.800 154.485 38.760 154.510 ;
        RECT 39.090 154.485 40.050 154.510 ;
        RECT 40.380 154.485 41.340 154.515 ;
        RECT 41.670 154.485 42.630 154.515 ;
        RECT 42.960 154.485 43.920 154.515 ;
        RECT 44.250 154.485 45.210 154.515 ;
        RECT 45.540 154.485 46.500 154.515 ;
        RECT 46.830 154.485 47.790 154.515 ;
        RECT 48.120 154.485 49.080 154.515 ;
        RECT 49.410 154.485 50.370 154.515 ;
        RECT 50.700 154.485 51.660 154.515 ;
        RECT 51.980 154.510 53.230 154.760 ;
        RECT 51.990 154.485 52.950 154.510 ;
        RECT 39.090 154.145 40.050 154.175 ;
        RECT 40.480 154.145 41.030 154.310 ;
        RECT 42.960 154.145 43.920 154.175 ;
        RECT 44.250 154.145 45.210 154.175 ;
        RECT 48.120 154.145 49.080 154.175 ;
        RECT 49.410 154.145 50.370 154.175 ;
        RECT 39.070 153.975 50.390 154.145 ;
        RECT 39.090 153.945 40.050 153.975 ;
        RECT 37.530 153.785 37.780 153.810 ;
        RECT 37.520 152.785 37.780 153.785 ;
        RECT 38.810 153.760 39.040 153.785 ;
        RECT 38.580 152.810 39.230 153.760 ;
        RECT 40.100 153.260 40.330 153.785 ;
        RECT 40.480 153.410 41.030 153.975 ;
        RECT 42.960 153.945 43.920 153.975 ;
        RECT 44.250 153.945 45.210 153.975 ;
        RECT 48.120 153.945 49.080 153.975 ;
        RECT 49.410 153.945 50.370 153.975 ;
        RECT 41.390 153.760 41.620 153.785 ;
        RECT 42.680 153.760 42.910 153.785 ;
        RECT 43.970 153.760 44.200 153.785 ;
        RECT 45.260 153.760 45.490 153.785 ;
        RECT 46.550 153.760 46.780 153.785 ;
        RECT 47.840 153.760 48.070 153.785 ;
        RECT 49.130 153.760 49.360 153.785 ;
        RECT 39.880 152.810 40.530 153.260 ;
        RECT 41.180 152.810 41.830 153.760 ;
        RECT 42.480 152.810 43.130 153.760 ;
        RECT 43.730 152.810 44.380 153.760 ;
        RECT 45.080 152.810 45.730 153.760 ;
        RECT 46.330 152.810 46.980 153.760 ;
        RECT 47.630 152.810 48.280 153.760 ;
        RECT 48.930 152.810 49.580 153.760 ;
        RECT 50.420 153.210 50.650 153.785 ;
        RECT 50.830 153.360 51.330 154.310 ;
        RECT 51.710 153.760 51.940 153.785 ;
        RECT 50.180 152.810 50.830 153.210 ;
        RECT 38.810 152.785 39.040 152.810 ;
        RECT 40.100 152.785 40.330 152.810 ;
        RECT 41.390 152.785 41.620 152.810 ;
        RECT 42.680 152.785 42.910 152.810 ;
        RECT 43.970 152.785 44.200 152.810 ;
        RECT 45.260 152.785 45.490 152.810 ;
        RECT 46.550 152.785 46.780 152.810 ;
        RECT 47.840 152.785 48.070 152.810 ;
        RECT 49.130 152.785 49.360 152.810 ;
        RECT 50.420 152.785 50.650 152.810 ;
        RECT 37.530 152.760 37.780 152.785 ;
        RECT 37.530 152.625 37.880 152.760 ;
        RECT 50.980 152.625 51.330 153.360 ;
        RECT 51.480 152.810 52.130 153.760 ;
        RECT 51.710 152.785 51.940 152.810 ;
        RECT 52.980 152.760 53.230 153.810 ;
        RECT 52.830 152.625 53.230 152.760 ;
        RECT 37.530 152.610 38.760 152.625 ;
        RECT 37.530 152.110 38.780 152.610 ;
        RECT 40.380 152.595 41.340 152.625 ;
        RECT 41.670 152.595 42.630 152.625 ;
        RECT 45.540 152.595 46.500 152.625 ;
        RECT 46.830 152.595 47.790 152.625 ;
        RECT 50.700 152.595 51.660 152.625 ;
        RECT 51.990 152.610 53.230 152.625 ;
        RECT 40.360 152.425 51.680 152.595 ;
        RECT 40.380 152.395 41.340 152.425 ;
        RECT 41.670 152.395 42.630 152.425 ;
        RECT 45.540 152.395 46.500 152.425 ;
        RECT 46.830 152.395 47.790 152.425 ;
        RECT 50.700 152.395 51.660 152.425 ;
        RECT 37.530 151.710 41.380 152.110 ;
        RECT 44.780 152.060 45.980 152.210 ;
        RECT 51.930 152.110 53.230 152.610 ;
        RECT 41.630 151.760 49.130 152.060 ;
        RECT 44.780 151.710 45.980 151.760 ;
        RECT 37.530 151.610 41.480 151.710 ;
        RECT 37.530 151.605 41.600 151.610 ;
        RECT 37.520 151.185 41.620 151.605 ;
        RECT 42.580 151.185 43.030 151.610 ;
        RECT 34.780 150.360 36.980 151.060 ;
        RECT 37.530 150.760 41.600 151.185 ;
        RECT 43.730 150.760 44.430 151.610 ;
        RECT 45.155 151.160 45.605 151.710 ;
        RECT 49.380 151.610 53.230 152.110 ;
        RECT 46.330 150.760 47.030 151.610 ;
        RECT 47.755 151.185 48.130 151.610 ;
        RECT 49.130 150.760 53.230 151.610 ;
        RECT 37.530 150.210 53.230 150.760 ;
        RECT 54.180 148.860 55.180 157.860 ;
        RECT 29.680 147.860 55.180 148.860 ;
        RECT 55.680 147.360 56.680 159.360 ;
        RECT 57.980 156.160 59.280 158.760 ;
        RECT 63.580 158.460 64.880 159.560 ;
        RECT 64.435 158.445 64.665 158.460 ;
        RECT 65.725 158.445 65.955 159.445 ;
        RECT 66.780 158.460 68.080 159.560 ;
        RECT 68.280 158.460 73.480 159.560 ;
        RECT 67.015 158.445 67.245 158.460 ;
        RECT 64.715 158.260 65.675 158.285 ;
        RECT 66.005 158.260 66.965 158.285 ;
        RECT 69.280 158.260 73.480 158.460 ;
        RECT 91.840 158.980 120.340 159.980 ;
        RECT 127.940 159.680 131.040 160.080 ;
        RECT 127.940 159.180 128.440 159.680 ;
        RECT 130.540 159.180 131.040 159.680 ;
        RECT 132.940 159.180 137.140 159.380 ;
        RECT 64.680 156.760 66.980 158.260 ;
        RECT 64.680 154.860 66.980 156.360 ;
        RECT 64.715 154.830 65.675 154.860 ;
        RECT 66.005 154.830 66.965 154.860 ;
        RECT 69.280 154.660 73.480 154.860 ;
        RECT 63.580 153.560 64.880 154.660 ;
        RECT 65.580 153.160 66.080 154.660 ;
        RECT 66.780 153.560 68.080 154.660 ;
        RECT 68.280 153.560 73.480 154.660 ;
        RECT 69.280 153.360 73.480 153.560 ;
        RECT 64.280 152.760 67.380 153.160 ;
        RECT 64.280 152.260 64.780 152.760 ;
        RECT 66.880 152.260 67.380 152.760 ;
        RECT 69.280 152.260 73.480 152.460 ;
        RECT 63.580 151.160 64.880 152.260 ;
        RECT 64.435 151.145 64.665 151.160 ;
        RECT 65.725 151.145 65.955 152.145 ;
        RECT 66.780 151.160 68.080 152.260 ;
        RECT 68.280 151.160 73.480 152.260 ;
        RECT 67.015 151.145 67.245 151.160 ;
        RECT 64.715 150.960 65.675 150.985 ;
        RECT 66.005 150.960 66.965 150.985 ;
        RECT 69.280 150.960 73.480 151.160 ;
        RECT 57.180 148.360 57.880 150.760 ;
        RECT 64.680 149.460 66.980 150.960 ;
        RECT 62.870 147.380 67.930 147.860 ;
        RECT 28.180 146.360 56.680 147.360 ;
        RECT 91.840 146.980 92.840 158.980 ;
        RECT 93.340 157.480 118.840 158.480 ;
        RECT 93.340 148.480 94.340 157.480 ;
        RECT 98.440 155.780 116.890 156.380 ;
        RECT 101.190 155.540 101.490 155.780 ;
        RECT 101.180 154.540 101.490 155.540 ;
        RECT 102.440 155.530 102.740 155.580 ;
        RECT 102.240 154.580 102.990 155.530 ;
        RECT 103.540 154.580 104.190 155.780 ;
        RECT 105.050 155.530 105.280 155.540 ;
        RECT 104.840 154.580 105.490 155.530 ;
        RECT 106.140 154.580 106.790 155.780 ;
        RECT 101.190 154.335 101.490 154.540 ;
        RECT 102.440 154.530 102.990 154.580 ;
        RECT 103.760 154.540 103.990 154.580 ;
        RECT 105.050 154.540 105.280 154.580 ;
        RECT 106.340 154.540 106.570 154.580 ;
        RECT 102.740 154.335 102.990 154.530 ;
        RECT 107.390 154.335 108.040 155.580 ;
        RECT 108.690 154.580 109.340 155.780 ;
        RECT 110.210 155.530 110.440 155.540 ;
        RECT 109.990 154.580 110.640 155.530 ;
        RECT 111.290 154.580 111.940 155.780 ;
        RECT 108.920 154.540 109.150 154.580 ;
        RECT 110.210 154.540 110.440 154.580 ;
        RECT 111.500 154.540 111.730 154.580 ;
        RECT 112.590 154.335 113.240 155.580 ;
        RECT 113.890 154.580 114.540 155.780 ;
        RECT 116.690 155.540 116.890 155.780 ;
        RECT 115.370 155.530 115.600 155.540 ;
        RECT 115.140 154.580 115.790 155.530 ;
        RECT 114.080 154.540 114.310 154.580 ;
        RECT 115.370 154.540 115.600 154.580 ;
        RECT 116.660 154.540 116.890 155.540 ;
        RECT 116.690 154.380 116.890 154.540 ;
        RECT 101.190 154.330 102.420 154.335 ;
        RECT 101.190 154.130 102.440 154.330 ;
        RECT 102.740 154.305 103.710 154.335 ;
        RECT 104.040 154.305 105.000 154.335 ;
        RECT 105.330 154.305 106.290 154.335 ;
        RECT 106.620 154.305 108.870 154.335 ;
        RECT 109.200 154.305 110.160 154.335 ;
        RECT 110.490 154.305 111.450 154.335 ;
        RECT 111.780 154.305 114.030 154.335 ;
        RECT 114.360 154.305 115.320 154.335 ;
        RECT 102.730 154.135 115.340 154.305 ;
        RECT 102.740 154.130 103.710 154.135 ;
        RECT 101.460 154.105 102.420 154.130 ;
        RECT 102.750 154.105 103.710 154.130 ;
        RECT 104.040 154.105 105.000 154.135 ;
        RECT 105.330 154.105 106.290 154.135 ;
        RECT 106.620 154.105 107.580 154.135 ;
        RECT 107.910 154.105 108.870 154.135 ;
        RECT 109.200 154.105 110.160 154.135 ;
        RECT 110.490 154.105 111.450 154.135 ;
        RECT 111.780 154.105 112.740 154.135 ;
        RECT 113.070 154.105 114.030 154.135 ;
        RECT 114.360 154.105 115.320 154.135 ;
        RECT 115.640 154.130 116.890 154.380 ;
        RECT 115.650 154.105 116.610 154.130 ;
        RECT 102.750 153.765 103.710 153.795 ;
        RECT 104.140 153.765 104.690 153.930 ;
        RECT 106.620 153.765 107.580 153.795 ;
        RECT 107.910 153.765 108.870 153.795 ;
        RECT 111.780 153.765 112.740 153.795 ;
        RECT 113.070 153.765 114.030 153.795 ;
        RECT 102.730 153.595 114.050 153.765 ;
        RECT 102.750 153.565 103.710 153.595 ;
        RECT 101.190 153.405 101.440 153.430 ;
        RECT 101.180 152.405 101.440 153.405 ;
        RECT 102.470 153.380 102.700 153.405 ;
        RECT 102.240 152.430 102.890 153.380 ;
        RECT 103.760 152.880 103.990 153.405 ;
        RECT 104.140 153.030 104.690 153.595 ;
        RECT 106.620 153.565 107.580 153.595 ;
        RECT 107.910 153.565 108.870 153.595 ;
        RECT 111.780 153.565 112.740 153.595 ;
        RECT 113.070 153.565 114.030 153.595 ;
        RECT 105.050 153.380 105.280 153.405 ;
        RECT 106.340 153.380 106.570 153.405 ;
        RECT 107.630 153.380 107.860 153.405 ;
        RECT 108.920 153.380 109.150 153.405 ;
        RECT 110.210 153.380 110.440 153.405 ;
        RECT 111.500 153.380 111.730 153.405 ;
        RECT 112.790 153.380 113.020 153.405 ;
        RECT 103.540 152.430 104.190 152.880 ;
        RECT 104.840 152.430 105.490 153.380 ;
        RECT 106.140 152.430 106.790 153.380 ;
        RECT 107.390 152.430 108.040 153.380 ;
        RECT 108.740 152.430 109.390 153.380 ;
        RECT 109.990 152.430 110.640 153.380 ;
        RECT 111.290 152.430 111.940 153.380 ;
        RECT 112.590 152.430 113.240 153.380 ;
        RECT 114.080 152.830 114.310 153.405 ;
        RECT 114.490 152.980 114.990 153.930 ;
        RECT 115.370 153.380 115.600 153.405 ;
        RECT 113.840 152.430 114.490 152.830 ;
        RECT 102.470 152.405 102.700 152.430 ;
        RECT 103.760 152.405 103.990 152.430 ;
        RECT 105.050 152.405 105.280 152.430 ;
        RECT 106.340 152.405 106.570 152.430 ;
        RECT 107.630 152.405 107.860 152.430 ;
        RECT 108.920 152.405 109.150 152.430 ;
        RECT 110.210 152.405 110.440 152.430 ;
        RECT 111.500 152.405 111.730 152.430 ;
        RECT 112.790 152.405 113.020 152.430 ;
        RECT 114.080 152.405 114.310 152.430 ;
        RECT 101.190 152.380 101.440 152.405 ;
        RECT 101.190 152.245 101.540 152.380 ;
        RECT 114.640 152.245 114.990 152.980 ;
        RECT 115.140 152.430 115.790 153.380 ;
        RECT 115.370 152.405 115.600 152.430 ;
        RECT 116.640 152.380 116.890 153.430 ;
        RECT 116.490 152.245 116.890 152.380 ;
        RECT 101.190 152.230 102.420 152.245 ;
        RECT 101.190 151.730 102.440 152.230 ;
        RECT 104.040 152.215 105.000 152.245 ;
        RECT 105.330 152.215 106.290 152.245 ;
        RECT 109.200 152.215 110.160 152.245 ;
        RECT 110.490 152.215 111.450 152.245 ;
        RECT 114.360 152.215 115.320 152.245 ;
        RECT 115.650 152.230 116.890 152.245 ;
        RECT 104.020 152.045 115.340 152.215 ;
        RECT 104.040 152.015 105.000 152.045 ;
        RECT 105.330 152.015 106.290 152.045 ;
        RECT 109.200 152.015 110.160 152.045 ;
        RECT 110.490 152.015 111.450 152.045 ;
        RECT 114.360 152.015 115.320 152.045 ;
        RECT 101.190 151.330 105.040 151.730 ;
        RECT 108.440 151.680 109.640 151.830 ;
        RECT 115.590 151.730 116.890 152.230 ;
        RECT 105.290 151.380 112.790 151.680 ;
        RECT 108.440 151.330 109.640 151.380 ;
        RECT 101.190 151.230 105.140 151.330 ;
        RECT 101.190 151.225 105.260 151.230 ;
        RECT 101.180 150.805 105.280 151.225 ;
        RECT 106.240 150.805 106.690 151.230 ;
        RECT 98.440 149.980 100.640 150.680 ;
        RECT 101.190 150.380 105.260 150.805 ;
        RECT 107.390 150.380 108.090 151.230 ;
        RECT 108.815 150.780 109.265 151.330 ;
        RECT 113.040 151.230 116.890 151.730 ;
        RECT 109.990 150.380 110.690 151.230 ;
        RECT 111.415 150.805 111.790 151.230 ;
        RECT 112.790 150.380 116.890 151.230 ;
        RECT 101.190 149.830 116.890 150.380 ;
        RECT 117.840 148.480 118.840 157.480 ;
        RECT 93.340 147.480 118.840 148.480 ;
        RECT 119.340 146.980 120.340 158.980 ;
        RECT 121.640 155.780 122.940 158.380 ;
        RECT 127.240 158.080 128.540 159.180 ;
        RECT 128.095 158.065 128.325 158.080 ;
        RECT 129.385 158.065 129.615 159.065 ;
        RECT 130.440 158.080 131.740 159.180 ;
        RECT 131.940 158.080 137.140 159.180 ;
        RECT 130.675 158.065 130.905 158.080 ;
        RECT 128.375 157.880 129.335 157.905 ;
        RECT 129.665 157.880 130.625 157.905 ;
        RECT 132.940 157.880 137.140 158.080 ;
        RECT 128.340 156.380 130.640 157.880 ;
        RECT 128.340 154.480 130.640 155.980 ;
        RECT 128.375 154.450 129.335 154.480 ;
        RECT 129.665 154.450 130.625 154.480 ;
        RECT 132.940 154.280 137.140 154.480 ;
        RECT 127.240 153.180 128.540 154.280 ;
        RECT 129.240 152.780 129.740 154.280 ;
        RECT 130.440 153.180 131.740 154.280 ;
        RECT 131.940 153.180 137.140 154.280 ;
        RECT 132.940 152.980 137.140 153.180 ;
        RECT 127.940 152.380 131.040 152.780 ;
        RECT 127.940 151.880 128.440 152.380 ;
        RECT 130.540 151.880 131.040 152.380 ;
        RECT 132.940 151.880 137.140 152.080 ;
        RECT 127.240 150.780 128.540 151.880 ;
        RECT 128.095 150.765 128.325 150.780 ;
        RECT 129.385 150.765 129.615 151.765 ;
        RECT 130.440 150.780 131.740 151.880 ;
        RECT 131.940 150.780 137.140 151.880 ;
        RECT 130.675 150.765 130.905 150.780 ;
        RECT 128.375 150.580 129.335 150.605 ;
        RECT 129.665 150.580 130.625 150.605 ;
        RECT 132.940 150.580 137.140 150.780 ;
        RECT 120.840 147.980 121.540 150.380 ;
        RECT 128.340 149.080 130.640 150.580 ;
        RECT 126.530 147.000 131.590 147.480 ;
        RECT 47.680 145.160 53.480 145.760 ;
        RECT 58.080 145.060 59.080 146.460 ;
        RECT 61.080 145.560 66.080 146.660 ;
        RECT 66.580 145.560 68.580 146.660 ;
        RECT 91.840 145.980 120.340 146.980 ;
        RECT 48.240 144.340 50.345 144.590 ;
        RECT 54.180 143.960 59.080 145.060 ;
        RECT 62.870 144.660 67.930 145.140 ;
        RECT 111.340 144.780 117.140 145.380 ;
        RECT 121.740 144.680 122.740 146.080 ;
        RECT 124.740 145.180 129.740 146.280 ;
        RECT 130.240 145.180 132.240 146.280 ;
        RECT 111.900 143.960 114.005 144.210 ;
        RECT 117.840 143.580 122.740 144.680 ;
        RECT 126.530 144.280 131.590 144.760 ;
        RECT 65.280 128.640 67.580 130.140 ;
        RECT 65.315 128.610 66.275 128.640 ;
        RECT 66.605 128.610 67.565 128.640 ;
        RECT 69.880 128.440 74.080 128.640 ;
        RECT 64.180 127.340 65.480 128.440 ;
        RECT 66.180 126.940 66.680 128.440 ;
        RECT 67.380 127.340 68.680 128.440 ;
        RECT 68.880 127.340 74.080 128.440 ;
        RECT 128.820 127.990 131.120 129.490 ;
        RECT 128.855 127.960 129.815 127.990 ;
        RECT 130.145 127.960 131.105 127.990 ;
        RECT 133.420 127.790 137.620 127.990 ;
        RECT 69.880 127.140 74.080 127.340 ;
        RECT 28.780 125.840 57.280 126.840 ;
        RECT 64.880 126.540 67.980 126.940 ;
        RECT 127.720 126.690 129.020 127.790 ;
        RECT 64.880 126.040 65.380 126.540 ;
        RECT 67.480 126.040 67.980 126.540 ;
        RECT 129.720 126.290 130.220 127.790 ;
        RECT 130.920 126.690 132.220 127.790 ;
        RECT 132.420 126.690 137.620 127.790 ;
        RECT 133.420 126.490 137.620 126.690 ;
        RECT 69.880 126.040 74.080 126.240 ;
        RECT 28.780 113.840 29.780 125.840 ;
        RECT 30.280 124.340 55.780 125.340 ;
        RECT 30.280 115.340 31.280 124.340 ;
        RECT 35.380 122.640 53.830 123.240 ;
        RECT 38.130 122.400 38.430 122.640 ;
        RECT 38.120 121.400 38.430 122.400 ;
        RECT 39.380 122.390 39.680 122.440 ;
        RECT 39.180 121.440 39.930 122.390 ;
        RECT 40.480 121.440 41.130 122.640 ;
        RECT 41.990 122.390 42.220 122.400 ;
        RECT 41.780 121.440 42.430 122.390 ;
        RECT 43.080 121.440 43.730 122.640 ;
        RECT 38.130 121.195 38.430 121.400 ;
        RECT 39.380 121.390 39.930 121.440 ;
        RECT 40.700 121.400 40.930 121.440 ;
        RECT 41.990 121.400 42.220 121.440 ;
        RECT 43.280 121.400 43.510 121.440 ;
        RECT 39.680 121.195 39.930 121.390 ;
        RECT 44.330 121.195 44.980 122.440 ;
        RECT 45.630 121.440 46.280 122.640 ;
        RECT 47.150 122.390 47.380 122.400 ;
        RECT 46.930 121.440 47.580 122.390 ;
        RECT 48.230 121.440 48.880 122.640 ;
        RECT 45.860 121.400 46.090 121.440 ;
        RECT 47.150 121.400 47.380 121.440 ;
        RECT 48.440 121.400 48.670 121.440 ;
        RECT 49.530 121.195 50.180 122.440 ;
        RECT 50.830 121.440 51.480 122.640 ;
        RECT 53.630 122.400 53.830 122.640 ;
        RECT 52.310 122.390 52.540 122.400 ;
        RECT 52.080 121.440 52.730 122.390 ;
        RECT 51.020 121.400 51.250 121.440 ;
        RECT 52.310 121.400 52.540 121.440 ;
        RECT 53.600 121.400 53.830 122.400 ;
        RECT 53.630 121.240 53.830 121.400 ;
        RECT 38.130 121.190 39.360 121.195 ;
        RECT 38.130 120.990 39.380 121.190 ;
        RECT 39.680 121.165 40.650 121.195 ;
        RECT 40.980 121.165 41.940 121.195 ;
        RECT 42.270 121.165 43.230 121.195 ;
        RECT 43.560 121.165 45.810 121.195 ;
        RECT 46.140 121.165 47.100 121.195 ;
        RECT 47.430 121.165 48.390 121.195 ;
        RECT 48.720 121.165 50.970 121.195 ;
        RECT 51.300 121.165 52.260 121.195 ;
        RECT 39.670 120.995 52.280 121.165 ;
        RECT 39.680 120.990 40.650 120.995 ;
        RECT 38.400 120.965 39.360 120.990 ;
        RECT 39.690 120.965 40.650 120.990 ;
        RECT 40.980 120.965 41.940 120.995 ;
        RECT 42.270 120.965 43.230 120.995 ;
        RECT 43.560 120.965 44.520 120.995 ;
        RECT 44.850 120.965 45.810 120.995 ;
        RECT 46.140 120.965 47.100 120.995 ;
        RECT 47.430 120.965 48.390 120.995 ;
        RECT 48.720 120.965 49.680 120.995 ;
        RECT 50.010 120.965 50.970 120.995 ;
        RECT 51.300 120.965 52.260 120.995 ;
        RECT 52.580 120.990 53.830 121.240 ;
        RECT 52.590 120.965 53.550 120.990 ;
        RECT 39.690 120.625 40.650 120.655 ;
        RECT 41.080 120.625 41.630 120.790 ;
        RECT 43.560 120.625 44.520 120.655 ;
        RECT 44.850 120.625 45.810 120.655 ;
        RECT 48.720 120.625 49.680 120.655 ;
        RECT 50.010 120.625 50.970 120.655 ;
        RECT 39.670 120.455 50.990 120.625 ;
        RECT 39.690 120.425 40.650 120.455 ;
        RECT 38.130 120.265 38.380 120.290 ;
        RECT 38.120 119.265 38.380 120.265 ;
        RECT 39.410 120.240 39.640 120.265 ;
        RECT 39.180 119.290 39.830 120.240 ;
        RECT 40.700 119.740 40.930 120.265 ;
        RECT 41.080 119.890 41.630 120.455 ;
        RECT 43.560 120.425 44.520 120.455 ;
        RECT 44.850 120.425 45.810 120.455 ;
        RECT 48.720 120.425 49.680 120.455 ;
        RECT 50.010 120.425 50.970 120.455 ;
        RECT 41.990 120.240 42.220 120.265 ;
        RECT 43.280 120.240 43.510 120.265 ;
        RECT 44.570 120.240 44.800 120.265 ;
        RECT 45.860 120.240 46.090 120.265 ;
        RECT 47.150 120.240 47.380 120.265 ;
        RECT 48.440 120.240 48.670 120.265 ;
        RECT 49.730 120.240 49.960 120.265 ;
        RECT 40.480 119.290 41.130 119.740 ;
        RECT 41.780 119.290 42.430 120.240 ;
        RECT 43.080 119.290 43.730 120.240 ;
        RECT 44.330 119.290 44.980 120.240 ;
        RECT 45.680 119.290 46.330 120.240 ;
        RECT 46.930 119.290 47.580 120.240 ;
        RECT 48.230 119.290 48.880 120.240 ;
        RECT 49.530 119.290 50.180 120.240 ;
        RECT 51.020 119.690 51.250 120.265 ;
        RECT 51.430 119.840 51.930 120.790 ;
        RECT 52.310 120.240 52.540 120.265 ;
        RECT 50.780 119.290 51.430 119.690 ;
        RECT 39.410 119.265 39.640 119.290 ;
        RECT 40.700 119.265 40.930 119.290 ;
        RECT 41.990 119.265 42.220 119.290 ;
        RECT 43.280 119.265 43.510 119.290 ;
        RECT 44.570 119.265 44.800 119.290 ;
        RECT 45.860 119.265 46.090 119.290 ;
        RECT 47.150 119.265 47.380 119.290 ;
        RECT 48.440 119.265 48.670 119.290 ;
        RECT 49.730 119.265 49.960 119.290 ;
        RECT 51.020 119.265 51.250 119.290 ;
        RECT 38.130 119.240 38.380 119.265 ;
        RECT 38.130 119.105 38.480 119.240 ;
        RECT 51.580 119.105 51.930 119.840 ;
        RECT 52.080 119.290 52.730 120.240 ;
        RECT 52.310 119.265 52.540 119.290 ;
        RECT 53.580 119.240 53.830 120.290 ;
        RECT 53.430 119.105 53.830 119.240 ;
        RECT 38.130 119.090 39.360 119.105 ;
        RECT 38.130 118.590 39.380 119.090 ;
        RECT 40.980 119.075 41.940 119.105 ;
        RECT 42.270 119.075 43.230 119.105 ;
        RECT 46.140 119.075 47.100 119.105 ;
        RECT 47.430 119.075 48.390 119.105 ;
        RECT 51.300 119.075 52.260 119.105 ;
        RECT 52.590 119.090 53.830 119.105 ;
        RECT 40.960 118.905 52.280 119.075 ;
        RECT 40.980 118.875 41.940 118.905 ;
        RECT 42.270 118.875 43.230 118.905 ;
        RECT 46.140 118.875 47.100 118.905 ;
        RECT 47.430 118.875 48.390 118.905 ;
        RECT 51.300 118.875 52.260 118.905 ;
        RECT 38.130 118.190 41.980 118.590 ;
        RECT 45.380 118.540 46.580 118.690 ;
        RECT 52.530 118.590 53.830 119.090 ;
        RECT 42.230 118.240 49.730 118.540 ;
        RECT 45.380 118.190 46.580 118.240 ;
        RECT 38.130 118.090 42.080 118.190 ;
        RECT 38.130 118.085 42.200 118.090 ;
        RECT 38.120 117.665 42.220 118.085 ;
        RECT 43.180 117.665 43.630 118.090 ;
        RECT 35.380 116.840 37.580 117.540 ;
        RECT 38.130 117.240 42.200 117.665 ;
        RECT 44.330 117.240 45.030 118.090 ;
        RECT 45.755 117.640 46.205 118.190 ;
        RECT 49.980 118.090 53.830 118.590 ;
        RECT 46.930 117.240 47.630 118.090 ;
        RECT 48.355 117.665 48.730 118.090 ;
        RECT 49.730 117.240 53.830 118.090 ;
        RECT 38.130 116.690 53.830 117.240 ;
        RECT 54.780 115.340 55.780 124.340 ;
        RECT 30.280 114.340 55.780 115.340 ;
        RECT 56.280 113.840 57.280 125.840 ;
        RECT 58.580 122.640 59.880 125.240 ;
        RECT 64.180 124.940 65.480 126.040 ;
        RECT 65.035 124.925 65.265 124.940 ;
        RECT 66.325 124.925 66.555 125.925 ;
        RECT 67.380 124.940 68.680 126.040 ;
        RECT 68.880 124.940 74.080 126.040 ;
        RECT 67.615 124.925 67.845 124.940 ;
        RECT 65.315 124.740 66.275 124.765 ;
        RECT 66.605 124.740 67.565 124.765 ;
        RECT 69.880 124.740 74.080 124.940 ;
        RECT 92.320 125.190 120.820 126.190 ;
        RECT 128.420 125.890 131.520 126.290 ;
        RECT 128.420 125.390 128.920 125.890 ;
        RECT 131.020 125.390 131.520 125.890 ;
        RECT 133.420 125.390 137.620 125.590 ;
        RECT 65.280 123.240 67.580 124.740 ;
        RECT 65.280 121.340 67.580 122.840 ;
        RECT 65.315 121.310 66.275 121.340 ;
        RECT 66.605 121.310 67.565 121.340 ;
        RECT 69.880 121.140 74.080 121.340 ;
        RECT 64.180 120.040 65.480 121.140 ;
        RECT 66.180 119.640 66.680 121.140 ;
        RECT 67.380 120.040 68.680 121.140 ;
        RECT 68.880 120.040 74.080 121.140 ;
        RECT 69.880 119.840 74.080 120.040 ;
        RECT 64.880 119.240 67.980 119.640 ;
        RECT 64.880 118.740 65.380 119.240 ;
        RECT 67.480 118.740 67.980 119.240 ;
        RECT 69.880 118.740 74.080 118.940 ;
        RECT 64.180 117.640 65.480 118.740 ;
        RECT 65.035 117.625 65.265 117.640 ;
        RECT 66.325 117.625 66.555 118.625 ;
        RECT 67.380 117.640 68.680 118.740 ;
        RECT 68.880 117.640 74.080 118.740 ;
        RECT 67.615 117.625 67.845 117.640 ;
        RECT 65.315 117.440 66.275 117.465 ;
        RECT 66.605 117.440 67.565 117.465 ;
        RECT 69.880 117.440 74.080 117.640 ;
        RECT 57.780 114.840 58.480 117.240 ;
        RECT 65.280 115.940 67.580 117.440 ;
        RECT 63.470 113.860 68.530 114.340 ;
        RECT 28.780 112.840 57.280 113.840 ;
        RECT 92.320 113.190 93.320 125.190 ;
        RECT 93.820 123.690 119.320 124.690 ;
        RECT 93.820 114.690 94.820 123.690 ;
        RECT 98.920 121.990 117.370 122.590 ;
        RECT 101.670 121.750 101.970 121.990 ;
        RECT 101.660 120.750 101.970 121.750 ;
        RECT 102.920 121.740 103.220 121.790 ;
        RECT 102.720 120.790 103.470 121.740 ;
        RECT 104.020 120.790 104.670 121.990 ;
        RECT 105.530 121.740 105.760 121.750 ;
        RECT 105.320 120.790 105.970 121.740 ;
        RECT 106.620 120.790 107.270 121.990 ;
        RECT 101.670 120.545 101.970 120.750 ;
        RECT 102.920 120.740 103.470 120.790 ;
        RECT 104.240 120.750 104.470 120.790 ;
        RECT 105.530 120.750 105.760 120.790 ;
        RECT 106.820 120.750 107.050 120.790 ;
        RECT 103.220 120.545 103.470 120.740 ;
        RECT 107.870 120.545 108.520 121.790 ;
        RECT 109.170 120.790 109.820 121.990 ;
        RECT 110.690 121.740 110.920 121.750 ;
        RECT 110.470 120.790 111.120 121.740 ;
        RECT 111.770 120.790 112.420 121.990 ;
        RECT 109.400 120.750 109.630 120.790 ;
        RECT 110.690 120.750 110.920 120.790 ;
        RECT 111.980 120.750 112.210 120.790 ;
        RECT 113.070 120.545 113.720 121.790 ;
        RECT 114.370 120.790 115.020 121.990 ;
        RECT 117.170 121.750 117.370 121.990 ;
        RECT 115.850 121.740 116.080 121.750 ;
        RECT 115.620 120.790 116.270 121.740 ;
        RECT 114.560 120.750 114.790 120.790 ;
        RECT 115.850 120.750 116.080 120.790 ;
        RECT 117.140 120.750 117.370 121.750 ;
        RECT 117.170 120.590 117.370 120.750 ;
        RECT 101.670 120.540 102.900 120.545 ;
        RECT 101.670 120.340 102.920 120.540 ;
        RECT 103.220 120.515 104.190 120.545 ;
        RECT 104.520 120.515 105.480 120.545 ;
        RECT 105.810 120.515 106.770 120.545 ;
        RECT 107.100 120.515 109.350 120.545 ;
        RECT 109.680 120.515 110.640 120.545 ;
        RECT 110.970 120.515 111.930 120.545 ;
        RECT 112.260 120.515 114.510 120.545 ;
        RECT 114.840 120.515 115.800 120.545 ;
        RECT 103.210 120.345 115.820 120.515 ;
        RECT 103.220 120.340 104.190 120.345 ;
        RECT 101.940 120.315 102.900 120.340 ;
        RECT 103.230 120.315 104.190 120.340 ;
        RECT 104.520 120.315 105.480 120.345 ;
        RECT 105.810 120.315 106.770 120.345 ;
        RECT 107.100 120.315 108.060 120.345 ;
        RECT 108.390 120.315 109.350 120.345 ;
        RECT 109.680 120.315 110.640 120.345 ;
        RECT 110.970 120.315 111.930 120.345 ;
        RECT 112.260 120.315 113.220 120.345 ;
        RECT 113.550 120.315 114.510 120.345 ;
        RECT 114.840 120.315 115.800 120.345 ;
        RECT 116.120 120.340 117.370 120.590 ;
        RECT 116.130 120.315 117.090 120.340 ;
        RECT 103.230 119.975 104.190 120.005 ;
        RECT 104.620 119.975 105.170 120.140 ;
        RECT 107.100 119.975 108.060 120.005 ;
        RECT 108.390 119.975 109.350 120.005 ;
        RECT 112.260 119.975 113.220 120.005 ;
        RECT 113.550 119.975 114.510 120.005 ;
        RECT 103.210 119.805 114.530 119.975 ;
        RECT 103.230 119.775 104.190 119.805 ;
        RECT 101.670 119.615 101.920 119.640 ;
        RECT 101.660 118.615 101.920 119.615 ;
        RECT 102.950 119.590 103.180 119.615 ;
        RECT 102.720 118.640 103.370 119.590 ;
        RECT 104.240 119.090 104.470 119.615 ;
        RECT 104.620 119.240 105.170 119.805 ;
        RECT 107.100 119.775 108.060 119.805 ;
        RECT 108.390 119.775 109.350 119.805 ;
        RECT 112.260 119.775 113.220 119.805 ;
        RECT 113.550 119.775 114.510 119.805 ;
        RECT 105.530 119.590 105.760 119.615 ;
        RECT 106.820 119.590 107.050 119.615 ;
        RECT 108.110 119.590 108.340 119.615 ;
        RECT 109.400 119.590 109.630 119.615 ;
        RECT 110.690 119.590 110.920 119.615 ;
        RECT 111.980 119.590 112.210 119.615 ;
        RECT 113.270 119.590 113.500 119.615 ;
        RECT 104.020 118.640 104.670 119.090 ;
        RECT 105.320 118.640 105.970 119.590 ;
        RECT 106.620 118.640 107.270 119.590 ;
        RECT 107.870 118.640 108.520 119.590 ;
        RECT 109.220 118.640 109.870 119.590 ;
        RECT 110.470 118.640 111.120 119.590 ;
        RECT 111.770 118.640 112.420 119.590 ;
        RECT 113.070 118.640 113.720 119.590 ;
        RECT 114.560 119.040 114.790 119.615 ;
        RECT 114.970 119.190 115.470 120.140 ;
        RECT 115.850 119.590 116.080 119.615 ;
        RECT 114.320 118.640 114.970 119.040 ;
        RECT 102.950 118.615 103.180 118.640 ;
        RECT 104.240 118.615 104.470 118.640 ;
        RECT 105.530 118.615 105.760 118.640 ;
        RECT 106.820 118.615 107.050 118.640 ;
        RECT 108.110 118.615 108.340 118.640 ;
        RECT 109.400 118.615 109.630 118.640 ;
        RECT 110.690 118.615 110.920 118.640 ;
        RECT 111.980 118.615 112.210 118.640 ;
        RECT 113.270 118.615 113.500 118.640 ;
        RECT 114.560 118.615 114.790 118.640 ;
        RECT 101.670 118.590 101.920 118.615 ;
        RECT 101.670 118.455 102.020 118.590 ;
        RECT 115.120 118.455 115.470 119.190 ;
        RECT 115.620 118.640 116.270 119.590 ;
        RECT 115.850 118.615 116.080 118.640 ;
        RECT 117.120 118.590 117.370 119.640 ;
        RECT 116.970 118.455 117.370 118.590 ;
        RECT 101.670 118.440 102.900 118.455 ;
        RECT 101.670 117.940 102.920 118.440 ;
        RECT 104.520 118.425 105.480 118.455 ;
        RECT 105.810 118.425 106.770 118.455 ;
        RECT 109.680 118.425 110.640 118.455 ;
        RECT 110.970 118.425 111.930 118.455 ;
        RECT 114.840 118.425 115.800 118.455 ;
        RECT 116.130 118.440 117.370 118.455 ;
        RECT 104.500 118.255 115.820 118.425 ;
        RECT 104.520 118.225 105.480 118.255 ;
        RECT 105.810 118.225 106.770 118.255 ;
        RECT 109.680 118.225 110.640 118.255 ;
        RECT 110.970 118.225 111.930 118.255 ;
        RECT 114.840 118.225 115.800 118.255 ;
        RECT 101.670 117.540 105.520 117.940 ;
        RECT 108.920 117.890 110.120 118.040 ;
        RECT 116.070 117.940 117.370 118.440 ;
        RECT 105.770 117.590 113.270 117.890 ;
        RECT 108.920 117.540 110.120 117.590 ;
        RECT 101.670 117.440 105.620 117.540 ;
        RECT 101.670 117.435 105.740 117.440 ;
        RECT 101.660 117.015 105.760 117.435 ;
        RECT 106.720 117.015 107.170 117.440 ;
        RECT 98.920 116.190 101.120 116.890 ;
        RECT 101.670 116.590 105.740 117.015 ;
        RECT 107.870 116.590 108.570 117.440 ;
        RECT 109.295 116.990 109.745 117.540 ;
        RECT 113.520 117.440 117.370 117.940 ;
        RECT 110.470 116.590 111.170 117.440 ;
        RECT 111.895 117.015 112.270 117.440 ;
        RECT 113.270 116.590 117.370 117.440 ;
        RECT 101.670 116.040 117.370 116.590 ;
        RECT 118.320 114.690 119.320 123.690 ;
        RECT 93.820 113.690 119.320 114.690 ;
        RECT 119.820 113.190 120.820 125.190 ;
        RECT 122.120 121.990 123.420 124.590 ;
        RECT 127.720 124.290 129.020 125.390 ;
        RECT 128.575 124.275 128.805 124.290 ;
        RECT 129.865 124.275 130.095 125.275 ;
        RECT 130.920 124.290 132.220 125.390 ;
        RECT 132.420 124.290 137.620 125.390 ;
        RECT 131.155 124.275 131.385 124.290 ;
        RECT 128.855 124.090 129.815 124.115 ;
        RECT 130.145 124.090 131.105 124.115 ;
        RECT 133.420 124.090 137.620 124.290 ;
        RECT 128.820 122.590 131.120 124.090 ;
        RECT 128.820 120.690 131.120 122.190 ;
        RECT 128.855 120.660 129.815 120.690 ;
        RECT 130.145 120.660 131.105 120.690 ;
        RECT 133.420 120.490 137.620 120.690 ;
        RECT 127.720 119.390 129.020 120.490 ;
        RECT 129.720 118.990 130.220 120.490 ;
        RECT 130.920 119.390 132.220 120.490 ;
        RECT 132.420 119.390 137.620 120.490 ;
        RECT 133.420 119.190 137.620 119.390 ;
        RECT 128.420 118.590 131.520 118.990 ;
        RECT 128.420 118.090 128.920 118.590 ;
        RECT 131.020 118.090 131.520 118.590 ;
        RECT 133.420 118.090 137.620 118.290 ;
        RECT 127.720 116.990 129.020 118.090 ;
        RECT 128.575 116.975 128.805 116.990 ;
        RECT 129.865 116.975 130.095 117.975 ;
        RECT 130.920 116.990 132.220 118.090 ;
        RECT 132.420 116.990 137.620 118.090 ;
        RECT 131.155 116.975 131.385 116.990 ;
        RECT 128.855 116.790 129.815 116.815 ;
        RECT 130.145 116.790 131.105 116.815 ;
        RECT 133.420 116.790 137.620 116.990 ;
        RECT 121.320 114.190 122.020 116.590 ;
        RECT 128.820 115.290 131.120 116.790 ;
        RECT 127.010 113.210 132.070 113.690 ;
        RECT 48.280 111.640 54.080 112.240 ;
        RECT 58.680 111.540 59.680 112.940 ;
        RECT 61.680 112.040 66.680 113.140 ;
        RECT 67.180 112.040 69.180 113.140 ;
        RECT 92.320 112.190 120.820 113.190 ;
        RECT 48.840 110.820 50.945 111.070 ;
        RECT 54.780 110.440 59.680 111.540 ;
        RECT 63.470 111.140 68.530 111.620 ;
        RECT 111.820 110.990 117.620 111.590 ;
        RECT 122.220 110.890 123.220 112.290 ;
        RECT 125.220 111.390 130.220 112.490 ;
        RECT 130.720 111.390 132.720 112.490 ;
        RECT 112.380 110.170 114.485 110.420 ;
        RECT 118.320 109.790 123.220 110.890 ;
        RECT 127.010 110.490 132.070 110.970 ;
        RECT 64.660 93.410 66.960 94.910 ;
        RECT 64.695 93.380 65.655 93.410 ;
        RECT 65.985 93.380 66.945 93.410 ;
        RECT 69.260 93.210 73.460 93.410 ;
        RECT 63.560 92.110 64.860 93.210 ;
        RECT 65.560 91.710 66.060 93.210 ;
        RECT 66.760 92.110 68.060 93.210 ;
        RECT 68.260 92.110 73.460 93.210 ;
        RECT 130.570 92.760 132.870 94.260 ;
        RECT 130.605 92.730 131.565 92.760 ;
        RECT 131.895 92.730 132.855 92.760 ;
        RECT 135.170 92.560 139.370 92.760 ;
        RECT 69.260 91.910 73.460 92.110 ;
        RECT 28.160 90.610 56.660 91.610 ;
        RECT 64.260 91.310 67.360 91.710 ;
        RECT 129.470 91.460 130.770 92.560 ;
        RECT 64.260 90.810 64.760 91.310 ;
        RECT 66.860 90.810 67.360 91.310 ;
        RECT 131.470 91.060 131.970 92.560 ;
        RECT 132.670 91.460 133.970 92.560 ;
        RECT 134.170 91.460 139.370 92.560 ;
        RECT 135.170 91.260 139.370 91.460 ;
        RECT 69.260 90.810 73.460 91.010 ;
        RECT 28.160 78.610 29.160 90.610 ;
        RECT 29.660 89.110 55.160 90.110 ;
        RECT 29.660 80.110 30.660 89.110 ;
        RECT 34.760 87.410 53.210 88.010 ;
        RECT 37.510 87.170 37.810 87.410 ;
        RECT 37.500 86.170 37.810 87.170 ;
        RECT 38.760 87.160 39.060 87.210 ;
        RECT 38.560 86.210 39.310 87.160 ;
        RECT 39.860 86.210 40.510 87.410 ;
        RECT 41.370 87.160 41.600 87.170 ;
        RECT 41.160 86.210 41.810 87.160 ;
        RECT 42.460 86.210 43.110 87.410 ;
        RECT 37.510 85.965 37.810 86.170 ;
        RECT 38.760 86.160 39.310 86.210 ;
        RECT 40.080 86.170 40.310 86.210 ;
        RECT 41.370 86.170 41.600 86.210 ;
        RECT 42.660 86.170 42.890 86.210 ;
        RECT 39.060 85.965 39.310 86.160 ;
        RECT 43.710 85.965 44.360 87.210 ;
        RECT 45.010 86.210 45.660 87.410 ;
        RECT 46.530 87.160 46.760 87.170 ;
        RECT 46.310 86.210 46.960 87.160 ;
        RECT 47.610 86.210 48.260 87.410 ;
        RECT 45.240 86.170 45.470 86.210 ;
        RECT 46.530 86.170 46.760 86.210 ;
        RECT 47.820 86.170 48.050 86.210 ;
        RECT 48.910 85.965 49.560 87.210 ;
        RECT 50.210 86.210 50.860 87.410 ;
        RECT 53.010 87.170 53.210 87.410 ;
        RECT 51.690 87.160 51.920 87.170 ;
        RECT 51.460 86.210 52.110 87.160 ;
        RECT 50.400 86.170 50.630 86.210 ;
        RECT 51.690 86.170 51.920 86.210 ;
        RECT 52.980 86.170 53.210 87.170 ;
        RECT 53.010 86.010 53.210 86.170 ;
        RECT 37.510 85.960 38.740 85.965 ;
        RECT 37.510 85.760 38.760 85.960 ;
        RECT 39.060 85.935 40.030 85.965 ;
        RECT 40.360 85.935 41.320 85.965 ;
        RECT 41.650 85.935 42.610 85.965 ;
        RECT 42.940 85.935 45.190 85.965 ;
        RECT 45.520 85.935 46.480 85.965 ;
        RECT 46.810 85.935 47.770 85.965 ;
        RECT 48.100 85.935 50.350 85.965 ;
        RECT 50.680 85.935 51.640 85.965 ;
        RECT 39.050 85.765 51.660 85.935 ;
        RECT 39.060 85.760 40.030 85.765 ;
        RECT 37.780 85.735 38.740 85.760 ;
        RECT 39.070 85.735 40.030 85.760 ;
        RECT 40.360 85.735 41.320 85.765 ;
        RECT 41.650 85.735 42.610 85.765 ;
        RECT 42.940 85.735 43.900 85.765 ;
        RECT 44.230 85.735 45.190 85.765 ;
        RECT 45.520 85.735 46.480 85.765 ;
        RECT 46.810 85.735 47.770 85.765 ;
        RECT 48.100 85.735 49.060 85.765 ;
        RECT 49.390 85.735 50.350 85.765 ;
        RECT 50.680 85.735 51.640 85.765 ;
        RECT 51.960 85.760 53.210 86.010 ;
        RECT 51.970 85.735 52.930 85.760 ;
        RECT 39.070 85.395 40.030 85.425 ;
        RECT 40.460 85.395 41.010 85.560 ;
        RECT 42.940 85.395 43.900 85.425 ;
        RECT 44.230 85.395 45.190 85.425 ;
        RECT 48.100 85.395 49.060 85.425 ;
        RECT 49.390 85.395 50.350 85.425 ;
        RECT 39.050 85.225 50.370 85.395 ;
        RECT 39.070 85.195 40.030 85.225 ;
        RECT 37.510 85.035 37.760 85.060 ;
        RECT 37.500 84.035 37.760 85.035 ;
        RECT 38.790 85.010 39.020 85.035 ;
        RECT 38.560 84.060 39.210 85.010 ;
        RECT 40.080 84.510 40.310 85.035 ;
        RECT 40.460 84.660 41.010 85.225 ;
        RECT 42.940 85.195 43.900 85.225 ;
        RECT 44.230 85.195 45.190 85.225 ;
        RECT 48.100 85.195 49.060 85.225 ;
        RECT 49.390 85.195 50.350 85.225 ;
        RECT 41.370 85.010 41.600 85.035 ;
        RECT 42.660 85.010 42.890 85.035 ;
        RECT 43.950 85.010 44.180 85.035 ;
        RECT 45.240 85.010 45.470 85.035 ;
        RECT 46.530 85.010 46.760 85.035 ;
        RECT 47.820 85.010 48.050 85.035 ;
        RECT 49.110 85.010 49.340 85.035 ;
        RECT 39.860 84.060 40.510 84.510 ;
        RECT 41.160 84.060 41.810 85.010 ;
        RECT 42.460 84.060 43.110 85.010 ;
        RECT 43.710 84.060 44.360 85.010 ;
        RECT 45.060 84.060 45.710 85.010 ;
        RECT 46.310 84.060 46.960 85.010 ;
        RECT 47.610 84.060 48.260 85.010 ;
        RECT 48.910 84.060 49.560 85.010 ;
        RECT 50.400 84.460 50.630 85.035 ;
        RECT 50.810 84.610 51.310 85.560 ;
        RECT 51.690 85.010 51.920 85.035 ;
        RECT 50.160 84.060 50.810 84.460 ;
        RECT 38.790 84.035 39.020 84.060 ;
        RECT 40.080 84.035 40.310 84.060 ;
        RECT 41.370 84.035 41.600 84.060 ;
        RECT 42.660 84.035 42.890 84.060 ;
        RECT 43.950 84.035 44.180 84.060 ;
        RECT 45.240 84.035 45.470 84.060 ;
        RECT 46.530 84.035 46.760 84.060 ;
        RECT 47.820 84.035 48.050 84.060 ;
        RECT 49.110 84.035 49.340 84.060 ;
        RECT 50.400 84.035 50.630 84.060 ;
        RECT 37.510 84.010 37.760 84.035 ;
        RECT 37.510 83.875 37.860 84.010 ;
        RECT 50.960 83.875 51.310 84.610 ;
        RECT 51.460 84.060 52.110 85.010 ;
        RECT 51.690 84.035 51.920 84.060 ;
        RECT 52.960 84.010 53.210 85.060 ;
        RECT 52.810 83.875 53.210 84.010 ;
        RECT 37.510 83.860 38.740 83.875 ;
        RECT 37.510 83.360 38.760 83.860 ;
        RECT 40.360 83.845 41.320 83.875 ;
        RECT 41.650 83.845 42.610 83.875 ;
        RECT 45.520 83.845 46.480 83.875 ;
        RECT 46.810 83.845 47.770 83.875 ;
        RECT 50.680 83.845 51.640 83.875 ;
        RECT 51.970 83.860 53.210 83.875 ;
        RECT 40.340 83.675 51.660 83.845 ;
        RECT 40.360 83.645 41.320 83.675 ;
        RECT 41.650 83.645 42.610 83.675 ;
        RECT 45.520 83.645 46.480 83.675 ;
        RECT 46.810 83.645 47.770 83.675 ;
        RECT 50.680 83.645 51.640 83.675 ;
        RECT 37.510 82.960 41.360 83.360 ;
        RECT 44.760 83.310 45.960 83.460 ;
        RECT 51.910 83.360 53.210 83.860 ;
        RECT 41.610 83.010 49.110 83.310 ;
        RECT 44.760 82.960 45.960 83.010 ;
        RECT 37.510 82.860 41.460 82.960 ;
        RECT 37.510 82.855 41.580 82.860 ;
        RECT 37.500 82.435 41.600 82.855 ;
        RECT 42.560 82.435 43.010 82.860 ;
        RECT 34.760 81.610 36.960 82.310 ;
        RECT 37.510 82.010 41.580 82.435 ;
        RECT 43.710 82.010 44.410 82.860 ;
        RECT 45.135 82.410 45.585 82.960 ;
        RECT 49.360 82.860 53.210 83.360 ;
        RECT 46.310 82.010 47.010 82.860 ;
        RECT 47.735 82.435 48.110 82.860 ;
        RECT 49.110 82.010 53.210 82.860 ;
        RECT 37.510 81.460 53.210 82.010 ;
        RECT 54.160 80.110 55.160 89.110 ;
        RECT 29.660 79.110 55.160 80.110 ;
        RECT 55.660 78.610 56.660 90.610 ;
        RECT 57.960 87.410 59.260 90.010 ;
        RECT 63.560 89.710 64.860 90.810 ;
        RECT 64.415 89.695 64.645 89.710 ;
        RECT 65.705 89.695 65.935 90.695 ;
        RECT 66.760 89.710 68.060 90.810 ;
        RECT 68.260 89.710 73.460 90.810 ;
        RECT 66.995 89.695 67.225 89.710 ;
        RECT 64.695 89.510 65.655 89.535 ;
        RECT 65.985 89.510 66.945 89.535 ;
        RECT 69.260 89.510 73.460 89.710 ;
        RECT 94.070 89.960 122.570 90.960 ;
        RECT 130.170 90.660 133.270 91.060 ;
        RECT 130.170 90.160 130.670 90.660 ;
        RECT 132.770 90.160 133.270 90.660 ;
        RECT 135.170 90.160 139.370 90.360 ;
        RECT 64.660 88.010 66.960 89.510 ;
        RECT 64.660 86.110 66.960 87.610 ;
        RECT 64.695 86.080 65.655 86.110 ;
        RECT 65.985 86.080 66.945 86.110 ;
        RECT 69.260 85.910 73.460 86.110 ;
        RECT 63.560 84.810 64.860 85.910 ;
        RECT 65.560 84.410 66.060 85.910 ;
        RECT 66.760 84.810 68.060 85.910 ;
        RECT 68.260 84.810 73.460 85.910 ;
        RECT 69.260 84.610 73.460 84.810 ;
        RECT 64.260 84.010 67.360 84.410 ;
        RECT 64.260 83.510 64.760 84.010 ;
        RECT 66.860 83.510 67.360 84.010 ;
        RECT 69.260 83.510 73.460 83.710 ;
        RECT 63.560 82.410 64.860 83.510 ;
        RECT 64.415 82.395 64.645 82.410 ;
        RECT 65.705 82.395 65.935 83.395 ;
        RECT 66.760 82.410 68.060 83.510 ;
        RECT 68.260 82.410 73.460 83.510 ;
        RECT 66.995 82.395 67.225 82.410 ;
        RECT 64.695 82.210 65.655 82.235 ;
        RECT 65.985 82.210 66.945 82.235 ;
        RECT 69.260 82.210 73.460 82.410 ;
        RECT 57.160 79.610 57.860 82.010 ;
        RECT 64.660 80.710 66.960 82.210 ;
        RECT 62.850 78.630 67.910 79.110 ;
        RECT 28.160 77.610 56.660 78.610 ;
        RECT 94.070 77.960 95.070 89.960 ;
        RECT 95.570 88.460 121.070 89.460 ;
        RECT 95.570 79.460 96.570 88.460 ;
        RECT 100.670 86.760 119.120 87.360 ;
        RECT 103.420 86.520 103.720 86.760 ;
        RECT 103.410 85.520 103.720 86.520 ;
        RECT 104.670 86.510 104.970 86.560 ;
        RECT 104.470 85.560 105.220 86.510 ;
        RECT 105.770 85.560 106.420 86.760 ;
        RECT 107.280 86.510 107.510 86.520 ;
        RECT 107.070 85.560 107.720 86.510 ;
        RECT 108.370 85.560 109.020 86.760 ;
        RECT 103.420 85.315 103.720 85.520 ;
        RECT 104.670 85.510 105.220 85.560 ;
        RECT 105.990 85.520 106.220 85.560 ;
        RECT 107.280 85.520 107.510 85.560 ;
        RECT 108.570 85.520 108.800 85.560 ;
        RECT 104.970 85.315 105.220 85.510 ;
        RECT 109.620 85.315 110.270 86.560 ;
        RECT 110.920 85.560 111.570 86.760 ;
        RECT 112.440 86.510 112.670 86.520 ;
        RECT 112.220 85.560 112.870 86.510 ;
        RECT 113.520 85.560 114.170 86.760 ;
        RECT 111.150 85.520 111.380 85.560 ;
        RECT 112.440 85.520 112.670 85.560 ;
        RECT 113.730 85.520 113.960 85.560 ;
        RECT 114.820 85.315 115.470 86.560 ;
        RECT 116.120 85.560 116.770 86.760 ;
        RECT 118.920 86.520 119.120 86.760 ;
        RECT 117.600 86.510 117.830 86.520 ;
        RECT 117.370 85.560 118.020 86.510 ;
        RECT 116.310 85.520 116.540 85.560 ;
        RECT 117.600 85.520 117.830 85.560 ;
        RECT 118.890 85.520 119.120 86.520 ;
        RECT 118.920 85.360 119.120 85.520 ;
        RECT 103.420 85.310 104.650 85.315 ;
        RECT 103.420 85.110 104.670 85.310 ;
        RECT 104.970 85.285 105.940 85.315 ;
        RECT 106.270 85.285 107.230 85.315 ;
        RECT 107.560 85.285 108.520 85.315 ;
        RECT 108.850 85.285 111.100 85.315 ;
        RECT 111.430 85.285 112.390 85.315 ;
        RECT 112.720 85.285 113.680 85.315 ;
        RECT 114.010 85.285 116.260 85.315 ;
        RECT 116.590 85.285 117.550 85.315 ;
        RECT 104.960 85.115 117.570 85.285 ;
        RECT 104.970 85.110 105.940 85.115 ;
        RECT 103.690 85.085 104.650 85.110 ;
        RECT 104.980 85.085 105.940 85.110 ;
        RECT 106.270 85.085 107.230 85.115 ;
        RECT 107.560 85.085 108.520 85.115 ;
        RECT 108.850 85.085 109.810 85.115 ;
        RECT 110.140 85.085 111.100 85.115 ;
        RECT 111.430 85.085 112.390 85.115 ;
        RECT 112.720 85.085 113.680 85.115 ;
        RECT 114.010 85.085 114.970 85.115 ;
        RECT 115.300 85.085 116.260 85.115 ;
        RECT 116.590 85.085 117.550 85.115 ;
        RECT 117.870 85.110 119.120 85.360 ;
        RECT 117.880 85.085 118.840 85.110 ;
        RECT 104.980 84.745 105.940 84.775 ;
        RECT 106.370 84.745 106.920 84.910 ;
        RECT 108.850 84.745 109.810 84.775 ;
        RECT 110.140 84.745 111.100 84.775 ;
        RECT 114.010 84.745 114.970 84.775 ;
        RECT 115.300 84.745 116.260 84.775 ;
        RECT 104.960 84.575 116.280 84.745 ;
        RECT 104.980 84.545 105.940 84.575 ;
        RECT 103.420 84.385 103.670 84.410 ;
        RECT 103.410 83.385 103.670 84.385 ;
        RECT 104.700 84.360 104.930 84.385 ;
        RECT 104.470 83.410 105.120 84.360 ;
        RECT 105.990 83.860 106.220 84.385 ;
        RECT 106.370 84.010 106.920 84.575 ;
        RECT 108.850 84.545 109.810 84.575 ;
        RECT 110.140 84.545 111.100 84.575 ;
        RECT 114.010 84.545 114.970 84.575 ;
        RECT 115.300 84.545 116.260 84.575 ;
        RECT 107.280 84.360 107.510 84.385 ;
        RECT 108.570 84.360 108.800 84.385 ;
        RECT 109.860 84.360 110.090 84.385 ;
        RECT 111.150 84.360 111.380 84.385 ;
        RECT 112.440 84.360 112.670 84.385 ;
        RECT 113.730 84.360 113.960 84.385 ;
        RECT 115.020 84.360 115.250 84.385 ;
        RECT 105.770 83.410 106.420 83.860 ;
        RECT 107.070 83.410 107.720 84.360 ;
        RECT 108.370 83.410 109.020 84.360 ;
        RECT 109.620 83.410 110.270 84.360 ;
        RECT 110.970 83.410 111.620 84.360 ;
        RECT 112.220 83.410 112.870 84.360 ;
        RECT 113.520 83.410 114.170 84.360 ;
        RECT 114.820 83.410 115.470 84.360 ;
        RECT 116.310 83.810 116.540 84.385 ;
        RECT 116.720 83.960 117.220 84.910 ;
        RECT 117.600 84.360 117.830 84.385 ;
        RECT 116.070 83.410 116.720 83.810 ;
        RECT 104.700 83.385 104.930 83.410 ;
        RECT 105.990 83.385 106.220 83.410 ;
        RECT 107.280 83.385 107.510 83.410 ;
        RECT 108.570 83.385 108.800 83.410 ;
        RECT 109.860 83.385 110.090 83.410 ;
        RECT 111.150 83.385 111.380 83.410 ;
        RECT 112.440 83.385 112.670 83.410 ;
        RECT 113.730 83.385 113.960 83.410 ;
        RECT 115.020 83.385 115.250 83.410 ;
        RECT 116.310 83.385 116.540 83.410 ;
        RECT 103.420 83.360 103.670 83.385 ;
        RECT 103.420 83.225 103.770 83.360 ;
        RECT 116.870 83.225 117.220 83.960 ;
        RECT 117.370 83.410 118.020 84.360 ;
        RECT 117.600 83.385 117.830 83.410 ;
        RECT 118.870 83.360 119.120 84.410 ;
        RECT 118.720 83.225 119.120 83.360 ;
        RECT 103.420 83.210 104.650 83.225 ;
        RECT 103.420 82.710 104.670 83.210 ;
        RECT 106.270 83.195 107.230 83.225 ;
        RECT 107.560 83.195 108.520 83.225 ;
        RECT 111.430 83.195 112.390 83.225 ;
        RECT 112.720 83.195 113.680 83.225 ;
        RECT 116.590 83.195 117.550 83.225 ;
        RECT 117.880 83.210 119.120 83.225 ;
        RECT 106.250 83.025 117.570 83.195 ;
        RECT 106.270 82.995 107.230 83.025 ;
        RECT 107.560 82.995 108.520 83.025 ;
        RECT 111.430 82.995 112.390 83.025 ;
        RECT 112.720 82.995 113.680 83.025 ;
        RECT 116.590 82.995 117.550 83.025 ;
        RECT 103.420 82.310 107.270 82.710 ;
        RECT 110.670 82.660 111.870 82.810 ;
        RECT 117.820 82.710 119.120 83.210 ;
        RECT 107.520 82.360 115.020 82.660 ;
        RECT 110.670 82.310 111.870 82.360 ;
        RECT 103.420 82.210 107.370 82.310 ;
        RECT 103.420 82.205 107.490 82.210 ;
        RECT 103.410 81.785 107.510 82.205 ;
        RECT 108.470 81.785 108.920 82.210 ;
        RECT 100.670 80.960 102.870 81.660 ;
        RECT 103.420 81.360 107.490 81.785 ;
        RECT 109.620 81.360 110.320 82.210 ;
        RECT 111.045 81.760 111.495 82.310 ;
        RECT 115.270 82.210 119.120 82.710 ;
        RECT 112.220 81.360 112.920 82.210 ;
        RECT 113.645 81.785 114.020 82.210 ;
        RECT 115.020 81.360 119.120 82.210 ;
        RECT 103.420 80.810 119.120 81.360 ;
        RECT 120.070 79.460 121.070 88.460 ;
        RECT 95.570 78.460 121.070 79.460 ;
        RECT 121.570 77.960 122.570 89.960 ;
        RECT 123.870 86.760 125.170 89.360 ;
        RECT 129.470 89.060 130.770 90.160 ;
        RECT 130.325 89.045 130.555 89.060 ;
        RECT 131.615 89.045 131.845 90.045 ;
        RECT 132.670 89.060 133.970 90.160 ;
        RECT 134.170 89.060 139.370 90.160 ;
        RECT 132.905 89.045 133.135 89.060 ;
        RECT 130.605 88.860 131.565 88.885 ;
        RECT 131.895 88.860 132.855 88.885 ;
        RECT 135.170 88.860 139.370 89.060 ;
        RECT 130.570 87.360 132.870 88.860 ;
        RECT 130.570 85.460 132.870 86.960 ;
        RECT 130.605 85.430 131.565 85.460 ;
        RECT 131.895 85.430 132.855 85.460 ;
        RECT 135.170 85.260 139.370 85.460 ;
        RECT 129.470 84.160 130.770 85.260 ;
        RECT 131.470 83.760 131.970 85.260 ;
        RECT 132.670 84.160 133.970 85.260 ;
        RECT 134.170 84.160 139.370 85.260 ;
        RECT 135.170 83.960 139.370 84.160 ;
        RECT 130.170 83.360 133.270 83.760 ;
        RECT 130.170 82.860 130.670 83.360 ;
        RECT 132.770 82.860 133.270 83.360 ;
        RECT 135.170 82.860 139.370 83.060 ;
        RECT 129.470 81.760 130.770 82.860 ;
        RECT 130.325 81.745 130.555 81.760 ;
        RECT 131.615 81.745 131.845 82.745 ;
        RECT 132.670 81.760 133.970 82.860 ;
        RECT 134.170 81.760 139.370 82.860 ;
        RECT 132.905 81.745 133.135 81.760 ;
        RECT 130.605 81.560 131.565 81.585 ;
        RECT 131.895 81.560 132.855 81.585 ;
        RECT 135.170 81.560 139.370 81.760 ;
        RECT 123.070 78.960 123.770 81.360 ;
        RECT 130.570 80.060 132.870 81.560 ;
        RECT 128.760 77.980 133.820 78.460 ;
        RECT 47.660 76.410 53.460 77.010 ;
        RECT 58.060 76.310 59.060 77.710 ;
        RECT 61.060 76.810 66.060 77.910 ;
        RECT 66.560 76.810 68.560 77.910 ;
        RECT 94.070 76.960 122.570 77.960 ;
        RECT 48.220 75.590 50.325 75.840 ;
        RECT 54.160 75.210 59.060 76.310 ;
        RECT 62.850 75.910 67.910 76.390 ;
        RECT 113.570 75.760 119.370 76.360 ;
        RECT 123.970 75.660 124.970 77.060 ;
        RECT 126.970 76.160 131.970 77.260 ;
        RECT 132.470 76.160 134.470 77.260 ;
        RECT 114.130 74.940 116.235 75.190 ;
        RECT 120.070 74.560 124.970 75.660 ;
        RECT 128.760 75.260 133.820 75.740 ;
      LAYER via ;
        RECT 64.550 192.100 66.650 193.000 ;
        RECT 128.620 192.880 130.720 193.780 ;
        RECT 63.450 190.400 64.550 191.300 ;
        RECT 66.650 190.400 67.750 191.300 ;
        RECT 72.650 190.200 73.050 191.300 ;
        RECT 127.520 191.180 128.620 192.080 ;
        RECT 130.720 191.180 131.820 192.080 ;
        RECT 136.720 190.980 137.120 192.080 ;
        RECT 37.100 188.900 53.150 189.700 ;
        RECT 101.170 189.680 117.220 190.480 ;
        RECT 37.100 185.700 52.900 186.100 ;
        RECT 38.400 184.450 38.950 184.750 ;
        RECT 41.000 184.450 41.550 184.750 ;
        RECT 43.550 184.200 44.100 184.750 ;
        RECT 46.150 184.450 46.700 184.800 ;
        RECT 48.750 184.200 49.300 184.800 ;
        RECT 51.300 184.450 51.850 184.800 ;
        RECT 38.400 182.850 38.950 183.150 ;
        RECT 40.300 182.900 40.750 183.700 ;
        RECT 41.000 182.850 41.550 183.150 ;
        RECT 39.700 182.300 40.250 182.600 ;
        RECT 42.300 182.300 42.850 182.600 ;
        RECT 43.550 182.850 44.100 183.150 ;
        RECT 44.900 182.300 45.450 182.600 ;
        RECT 46.150 182.850 46.700 183.150 ;
        RECT 47.450 182.300 48.000 182.600 ;
        RECT 48.750 182.850 49.300 183.150 ;
        RECT 50.650 182.950 51.050 183.700 ;
        RECT 50.000 182.300 50.550 182.600 ;
        RECT 51.300 182.850 51.850 183.150 ;
        RECT 44.600 181.350 45.700 181.650 ;
        RECT 42.425 180.675 42.700 181.050 ;
        RECT 34.600 179.850 36.700 180.450 ;
        RECT 47.575 180.675 47.850 181.050 ;
        RECT 37.400 179.750 52.900 180.100 ;
        RECT 37.100 177.400 53.150 178.200 ;
        RECT 57.850 185.700 58.950 188.100 ;
        RECT 63.450 188.000 64.550 188.900 ;
        RECT 66.650 188.000 67.750 188.900 ;
        RECT 71.750 187.900 72.150 189.000 ;
        RECT 64.550 186.300 66.650 187.200 ;
        RECT 64.550 184.800 66.650 185.700 ;
        RECT 63.450 183.100 64.550 184.000 ;
        RECT 66.650 183.100 67.750 184.000 ;
        RECT 72.650 182.900 73.050 184.000 ;
        RECT 63.450 180.700 64.550 181.600 ;
        RECT 66.650 180.700 67.750 181.600 ;
        RECT 71.750 180.600 72.150 181.700 ;
        RECT 57.050 177.900 57.550 180.100 ;
        RECT 64.550 179.000 66.650 179.900 ;
        RECT 101.170 186.480 116.970 186.880 ;
        RECT 102.470 185.230 103.020 185.530 ;
        RECT 105.070 185.230 105.620 185.530 ;
        RECT 107.620 184.980 108.170 185.530 ;
        RECT 110.220 185.230 110.770 185.580 ;
        RECT 112.820 184.980 113.370 185.580 ;
        RECT 115.370 185.230 115.920 185.580 ;
        RECT 102.470 183.630 103.020 183.930 ;
        RECT 104.370 183.680 104.820 184.480 ;
        RECT 105.070 183.630 105.620 183.930 ;
        RECT 103.770 183.080 104.320 183.380 ;
        RECT 106.370 183.080 106.920 183.380 ;
        RECT 107.620 183.630 108.170 183.930 ;
        RECT 108.970 183.080 109.520 183.380 ;
        RECT 110.220 183.630 110.770 183.930 ;
        RECT 111.520 183.080 112.070 183.380 ;
        RECT 112.820 183.630 113.370 183.930 ;
        RECT 114.720 183.730 115.120 184.480 ;
        RECT 114.070 183.080 114.620 183.380 ;
        RECT 115.370 183.630 115.920 183.930 ;
        RECT 108.670 182.130 109.770 182.430 ;
        RECT 106.495 181.455 106.770 181.830 ;
        RECT 98.670 180.630 100.770 181.230 ;
        RECT 111.645 181.455 111.920 181.830 ;
        RECT 101.470 180.530 116.970 180.880 ;
        RECT 101.170 178.180 117.220 178.980 ;
        RECT 121.920 186.480 123.020 188.880 ;
        RECT 127.520 188.780 128.620 189.680 ;
        RECT 130.720 188.780 131.820 189.680 ;
        RECT 135.820 188.680 136.220 189.780 ;
        RECT 128.620 187.080 130.720 187.980 ;
        RECT 128.620 185.580 130.720 186.480 ;
        RECT 127.520 183.880 128.620 184.780 ;
        RECT 130.720 183.880 131.820 184.780 ;
        RECT 136.720 183.680 137.120 184.780 ;
        RECT 127.520 181.480 128.620 182.380 ;
        RECT 130.720 181.480 131.820 182.380 ;
        RECT 135.820 181.380 136.220 182.480 ;
        RECT 121.120 178.680 121.620 180.880 ;
        RECT 128.620 179.780 130.720 180.680 ;
        RECT 126.820 177.680 131.620 177.980 ;
        RECT 62.750 176.900 67.550 177.200 ;
        RECT 47.550 174.700 53.150 175.100 ;
        RECT 57.950 174.400 58.750 175.800 ;
        RECT 54.050 173.500 58.750 174.400 ;
        RECT 60.950 175.100 61.850 176.000 ;
        RECT 67.350 175.100 68.250 176.000 ;
        RECT 111.620 175.480 117.220 175.880 ;
        RECT 122.020 175.180 122.820 176.580 ;
        RECT 62.750 174.200 67.650 174.500 ;
        RECT 118.120 174.280 122.820 175.180 ;
        RECT 125.020 175.880 125.920 176.780 ;
        RECT 131.420 175.880 132.320 176.780 ;
        RECT 126.820 174.980 131.720 175.280 ;
        RECT 64.780 162.660 66.880 163.560 ;
        RECT 128.440 162.280 130.540 163.180 ;
        RECT 63.680 160.960 64.780 161.860 ;
        RECT 66.880 160.960 67.980 161.860 ;
        RECT 72.880 160.760 73.280 161.860 ;
        RECT 127.340 160.580 128.440 161.480 ;
        RECT 37.330 159.460 53.380 160.260 ;
        RECT 130.540 160.580 131.640 161.480 ;
        RECT 136.540 160.380 136.940 161.480 ;
        RECT 37.330 156.260 53.130 156.660 ;
        RECT 38.630 155.010 39.180 155.310 ;
        RECT 41.230 155.010 41.780 155.310 ;
        RECT 43.780 154.760 44.330 155.310 ;
        RECT 46.380 155.010 46.930 155.360 ;
        RECT 48.980 154.760 49.530 155.360 ;
        RECT 51.530 155.010 52.080 155.360 ;
        RECT 38.630 153.410 39.180 153.710 ;
        RECT 40.530 153.460 40.980 154.260 ;
        RECT 41.230 153.410 41.780 153.710 ;
        RECT 39.930 152.860 40.480 153.160 ;
        RECT 42.530 152.860 43.080 153.160 ;
        RECT 43.780 153.410 44.330 153.710 ;
        RECT 45.130 152.860 45.680 153.160 ;
        RECT 46.380 153.410 46.930 153.710 ;
        RECT 47.680 152.860 48.230 153.160 ;
        RECT 48.980 153.410 49.530 153.710 ;
        RECT 50.880 153.510 51.280 154.260 ;
        RECT 50.230 152.860 50.780 153.160 ;
        RECT 51.530 153.410 52.080 153.710 ;
        RECT 44.830 151.910 45.930 152.210 ;
        RECT 42.655 151.235 42.930 151.610 ;
        RECT 34.830 150.410 36.930 151.010 ;
        RECT 47.805 151.235 48.080 151.610 ;
        RECT 37.630 150.310 53.130 150.660 ;
        RECT 37.330 147.960 53.380 148.760 ;
        RECT 58.080 156.260 59.180 158.660 ;
        RECT 63.680 158.560 64.780 159.460 ;
        RECT 66.880 158.560 67.980 159.460 ;
        RECT 71.980 158.460 72.380 159.560 ;
        RECT 100.990 159.080 117.040 159.880 ;
        RECT 64.780 156.860 66.880 157.760 ;
        RECT 64.780 155.360 66.880 156.260 ;
        RECT 63.680 153.660 64.780 154.560 ;
        RECT 66.880 153.660 67.980 154.560 ;
        RECT 72.880 153.460 73.280 154.560 ;
        RECT 63.680 151.260 64.780 152.160 ;
        RECT 66.880 151.260 67.980 152.160 ;
        RECT 71.980 151.160 72.380 152.260 ;
        RECT 57.280 148.460 57.780 150.660 ;
        RECT 64.780 149.560 66.880 150.460 ;
        RECT 62.980 147.460 67.780 147.760 ;
        RECT 100.990 155.880 116.790 156.280 ;
        RECT 102.290 154.630 102.840 154.930 ;
        RECT 104.890 154.630 105.440 154.930 ;
        RECT 107.440 154.380 107.990 154.930 ;
        RECT 110.040 154.630 110.590 154.980 ;
        RECT 112.640 154.380 113.190 154.980 ;
        RECT 115.190 154.630 115.740 154.980 ;
        RECT 102.290 153.030 102.840 153.330 ;
        RECT 104.190 153.080 104.640 153.880 ;
        RECT 104.890 153.030 105.440 153.330 ;
        RECT 103.590 152.480 104.140 152.780 ;
        RECT 106.190 152.480 106.740 152.780 ;
        RECT 107.440 153.030 107.990 153.330 ;
        RECT 108.790 152.480 109.340 152.780 ;
        RECT 110.040 153.030 110.590 153.330 ;
        RECT 111.340 152.480 111.890 152.780 ;
        RECT 112.640 153.030 113.190 153.330 ;
        RECT 114.540 153.130 114.940 153.880 ;
        RECT 113.890 152.480 114.440 152.780 ;
        RECT 115.190 153.030 115.740 153.330 ;
        RECT 108.490 151.530 109.590 151.830 ;
        RECT 106.315 150.855 106.590 151.230 ;
        RECT 98.490 150.030 100.590 150.630 ;
        RECT 111.465 150.855 111.740 151.230 ;
        RECT 101.290 149.930 116.790 150.280 ;
        RECT 100.990 147.580 117.040 148.380 ;
        RECT 121.740 155.880 122.840 158.280 ;
        RECT 127.340 158.180 128.440 159.080 ;
        RECT 130.540 158.180 131.640 159.080 ;
        RECT 135.640 158.080 136.040 159.180 ;
        RECT 128.440 156.480 130.540 157.380 ;
        RECT 128.440 154.980 130.540 155.880 ;
        RECT 127.340 153.280 128.440 154.180 ;
        RECT 130.540 153.280 131.640 154.180 ;
        RECT 136.540 153.080 136.940 154.180 ;
        RECT 127.340 150.880 128.440 151.780 ;
        RECT 130.540 150.880 131.640 151.780 ;
        RECT 135.640 150.780 136.040 151.880 ;
        RECT 120.940 148.080 121.440 150.280 ;
        RECT 128.440 149.180 130.540 150.080 ;
        RECT 126.640 147.080 131.440 147.380 ;
        RECT 47.780 145.260 53.380 145.660 ;
        RECT 58.180 144.960 58.980 146.360 ;
        RECT 54.280 144.060 58.980 144.960 ;
        RECT 61.180 145.660 62.080 146.560 ;
        RECT 67.580 145.660 68.480 146.560 ;
        RECT 62.980 144.760 67.880 145.060 ;
        RECT 111.440 144.880 117.040 145.280 ;
        RECT 121.840 144.580 122.640 145.980 ;
        RECT 117.940 143.680 122.640 144.580 ;
        RECT 124.840 145.280 125.740 146.180 ;
        RECT 131.240 145.280 132.140 146.180 ;
        RECT 126.640 144.380 131.540 144.680 ;
        RECT 65.380 129.140 67.480 130.040 ;
        RECT 64.280 127.440 65.380 128.340 ;
        RECT 67.480 127.440 68.580 128.340 ;
        RECT 73.480 127.240 73.880 128.340 ;
        RECT 128.920 128.490 131.020 129.390 ;
        RECT 37.930 125.940 53.980 126.740 ;
        RECT 127.820 126.790 128.920 127.690 ;
        RECT 131.020 126.790 132.120 127.690 ;
        RECT 137.020 126.590 137.420 127.690 ;
        RECT 37.930 122.740 53.730 123.140 ;
        RECT 39.230 121.490 39.780 121.790 ;
        RECT 41.830 121.490 42.380 121.790 ;
        RECT 44.380 121.240 44.930 121.790 ;
        RECT 46.980 121.490 47.530 121.840 ;
        RECT 49.580 121.240 50.130 121.840 ;
        RECT 52.130 121.490 52.680 121.840 ;
        RECT 39.230 119.890 39.780 120.190 ;
        RECT 41.130 119.940 41.580 120.740 ;
        RECT 41.830 119.890 42.380 120.190 ;
        RECT 40.530 119.340 41.080 119.640 ;
        RECT 43.130 119.340 43.680 119.640 ;
        RECT 44.380 119.890 44.930 120.190 ;
        RECT 45.730 119.340 46.280 119.640 ;
        RECT 46.980 119.890 47.530 120.190 ;
        RECT 48.280 119.340 48.830 119.640 ;
        RECT 49.580 119.890 50.130 120.190 ;
        RECT 51.480 119.990 51.880 120.740 ;
        RECT 50.830 119.340 51.380 119.640 ;
        RECT 52.130 119.890 52.680 120.190 ;
        RECT 45.430 118.390 46.530 118.690 ;
        RECT 43.255 117.715 43.530 118.090 ;
        RECT 35.430 116.890 37.530 117.490 ;
        RECT 48.405 117.715 48.680 118.090 ;
        RECT 38.230 116.790 53.730 117.140 ;
        RECT 37.930 114.440 53.980 115.240 ;
        RECT 58.680 122.740 59.780 125.140 ;
        RECT 64.280 125.040 65.380 125.940 ;
        RECT 67.480 125.040 68.580 125.940 ;
        RECT 72.580 124.940 72.980 126.040 ;
        RECT 101.470 125.290 117.520 126.090 ;
        RECT 65.380 123.340 67.480 124.240 ;
        RECT 65.380 121.840 67.480 122.740 ;
        RECT 64.280 120.140 65.380 121.040 ;
        RECT 67.480 120.140 68.580 121.040 ;
        RECT 73.480 119.940 73.880 121.040 ;
        RECT 64.280 117.740 65.380 118.640 ;
        RECT 67.480 117.740 68.580 118.640 ;
        RECT 72.580 117.640 72.980 118.740 ;
        RECT 57.880 114.940 58.380 117.140 ;
        RECT 65.380 116.040 67.480 116.940 ;
        RECT 63.580 113.940 68.380 114.240 ;
        RECT 101.470 122.090 117.270 122.490 ;
        RECT 102.770 120.840 103.320 121.140 ;
        RECT 105.370 120.840 105.920 121.140 ;
        RECT 107.920 120.590 108.470 121.140 ;
        RECT 110.520 120.840 111.070 121.190 ;
        RECT 113.120 120.590 113.670 121.190 ;
        RECT 115.670 120.840 116.220 121.190 ;
        RECT 102.770 119.240 103.320 119.540 ;
        RECT 104.670 119.290 105.120 120.090 ;
        RECT 105.370 119.240 105.920 119.540 ;
        RECT 104.070 118.690 104.620 118.990 ;
        RECT 106.670 118.690 107.220 118.990 ;
        RECT 107.920 119.240 108.470 119.540 ;
        RECT 109.270 118.690 109.820 118.990 ;
        RECT 110.520 119.240 111.070 119.540 ;
        RECT 111.820 118.690 112.370 118.990 ;
        RECT 113.120 119.240 113.670 119.540 ;
        RECT 115.020 119.340 115.420 120.090 ;
        RECT 114.370 118.690 114.920 118.990 ;
        RECT 115.670 119.240 116.220 119.540 ;
        RECT 108.970 117.740 110.070 118.040 ;
        RECT 106.795 117.065 107.070 117.440 ;
        RECT 98.970 116.240 101.070 116.840 ;
        RECT 111.945 117.065 112.220 117.440 ;
        RECT 101.770 116.140 117.270 116.490 ;
        RECT 101.470 113.790 117.520 114.590 ;
        RECT 122.220 122.090 123.320 124.490 ;
        RECT 127.820 124.390 128.920 125.290 ;
        RECT 131.020 124.390 132.120 125.290 ;
        RECT 136.120 124.290 136.520 125.390 ;
        RECT 128.920 122.690 131.020 123.590 ;
        RECT 128.920 121.190 131.020 122.090 ;
        RECT 127.820 119.490 128.920 120.390 ;
        RECT 131.020 119.490 132.120 120.390 ;
        RECT 137.020 119.290 137.420 120.390 ;
        RECT 127.820 117.090 128.920 117.990 ;
        RECT 131.020 117.090 132.120 117.990 ;
        RECT 136.120 116.990 136.520 118.090 ;
        RECT 121.420 114.290 121.920 116.490 ;
        RECT 128.920 115.390 131.020 116.290 ;
        RECT 127.120 113.290 131.920 113.590 ;
        RECT 48.380 111.740 53.980 112.140 ;
        RECT 58.780 111.440 59.580 112.840 ;
        RECT 54.880 110.540 59.580 111.440 ;
        RECT 61.780 112.140 62.680 113.040 ;
        RECT 68.180 112.140 69.080 113.040 ;
        RECT 63.580 111.240 68.480 111.540 ;
        RECT 111.920 111.090 117.520 111.490 ;
        RECT 122.320 110.790 123.120 112.190 ;
        RECT 118.420 109.890 123.120 110.790 ;
        RECT 125.320 111.490 126.220 112.390 ;
        RECT 131.720 111.490 132.620 112.390 ;
        RECT 127.120 110.590 132.020 110.890 ;
        RECT 64.760 93.910 66.860 94.810 ;
        RECT 63.660 92.210 64.760 93.110 ;
        RECT 66.860 92.210 67.960 93.110 ;
        RECT 72.860 92.010 73.260 93.110 ;
        RECT 130.670 93.260 132.770 94.160 ;
        RECT 37.310 90.710 53.360 91.510 ;
        RECT 129.570 91.560 130.670 92.460 ;
        RECT 132.770 91.560 133.870 92.460 ;
        RECT 138.770 91.360 139.170 92.460 ;
        RECT 37.310 87.510 53.110 87.910 ;
        RECT 38.610 86.260 39.160 86.560 ;
        RECT 41.210 86.260 41.760 86.560 ;
        RECT 43.760 86.010 44.310 86.560 ;
        RECT 46.360 86.260 46.910 86.610 ;
        RECT 48.960 86.010 49.510 86.610 ;
        RECT 51.510 86.260 52.060 86.610 ;
        RECT 38.610 84.660 39.160 84.960 ;
        RECT 40.510 84.710 40.960 85.510 ;
        RECT 41.210 84.660 41.760 84.960 ;
        RECT 39.910 84.110 40.460 84.410 ;
        RECT 42.510 84.110 43.060 84.410 ;
        RECT 43.760 84.660 44.310 84.960 ;
        RECT 45.110 84.110 45.660 84.410 ;
        RECT 46.360 84.660 46.910 84.960 ;
        RECT 47.660 84.110 48.210 84.410 ;
        RECT 48.960 84.660 49.510 84.960 ;
        RECT 50.860 84.760 51.260 85.510 ;
        RECT 50.210 84.110 50.760 84.410 ;
        RECT 51.510 84.660 52.060 84.960 ;
        RECT 44.810 83.160 45.910 83.460 ;
        RECT 42.635 82.485 42.910 82.860 ;
        RECT 34.810 81.660 36.910 82.260 ;
        RECT 47.785 82.485 48.060 82.860 ;
        RECT 37.610 81.560 53.110 81.910 ;
        RECT 37.310 79.210 53.360 80.010 ;
        RECT 58.060 87.510 59.160 89.910 ;
        RECT 63.660 89.810 64.760 90.710 ;
        RECT 66.860 89.810 67.960 90.710 ;
        RECT 71.960 89.710 72.360 90.810 ;
        RECT 103.220 90.060 119.270 90.860 ;
        RECT 64.760 88.110 66.860 89.010 ;
        RECT 64.760 86.610 66.860 87.510 ;
        RECT 63.660 84.910 64.760 85.810 ;
        RECT 66.860 84.910 67.960 85.810 ;
        RECT 72.860 84.710 73.260 85.810 ;
        RECT 63.660 82.510 64.760 83.410 ;
        RECT 66.860 82.510 67.960 83.410 ;
        RECT 71.960 82.410 72.360 83.510 ;
        RECT 57.260 79.710 57.760 81.910 ;
        RECT 64.760 80.810 66.860 81.710 ;
        RECT 62.960 78.710 67.760 79.010 ;
        RECT 103.220 86.860 119.020 87.260 ;
        RECT 104.520 85.610 105.070 85.910 ;
        RECT 107.120 85.610 107.670 85.910 ;
        RECT 109.670 85.360 110.220 85.910 ;
        RECT 112.270 85.610 112.820 85.960 ;
        RECT 114.870 85.360 115.420 85.960 ;
        RECT 117.420 85.610 117.970 85.960 ;
        RECT 104.520 84.010 105.070 84.310 ;
        RECT 106.420 84.060 106.870 84.860 ;
        RECT 107.120 84.010 107.670 84.310 ;
        RECT 105.820 83.460 106.370 83.760 ;
        RECT 108.420 83.460 108.970 83.760 ;
        RECT 109.670 84.010 110.220 84.310 ;
        RECT 111.020 83.460 111.570 83.760 ;
        RECT 112.270 84.010 112.820 84.310 ;
        RECT 113.570 83.460 114.120 83.760 ;
        RECT 114.870 84.010 115.420 84.310 ;
        RECT 116.770 84.110 117.170 84.860 ;
        RECT 116.120 83.460 116.670 83.760 ;
        RECT 117.420 84.010 117.970 84.310 ;
        RECT 110.720 82.510 111.820 82.810 ;
        RECT 108.545 81.835 108.820 82.210 ;
        RECT 100.720 81.010 102.820 81.610 ;
        RECT 113.695 81.835 113.970 82.210 ;
        RECT 103.520 80.910 119.020 81.260 ;
        RECT 103.220 78.560 119.270 79.360 ;
        RECT 123.970 86.860 125.070 89.260 ;
        RECT 129.570 89.160 130.670 90.060 ;
        RECT 132.770 89.160 133.870 90.060 ;
        RECT 137.870 89.060 138.270 90.160 ;
        RECT 130.670 87.460 132.770 88.360 ;
        RECT 130.670 85.960 132.770 86.860 ;
        RECT 129.570 84.260 130.670 85.160 ;
        RECT 132.770 84.260 133.870 85.160 ;
        RECT 138.770 84.060 139.170 85.160 ;
        RECT 129.570 81.860 130.670 82.760 ;
        RECT 132.770 81.860 133.870 82.760 ;
        RECT 137.870 81.760 138.270 82.860 ;
        RECT 123.170 79.060 123.670 81.260 ;
        RECT 130.670 80.160 132.770 81.060 ;
        RECT 128.870 78.060 133.670 78.360 ;
        RECT 47.760 76.510 53.360 76.910 ;
        RECT 58.160 76.210 58.960 77.610 ;
        RECT 54.260 75.310 58.960 76.210 ;
        RECT 61.160 76.910 62.060 77.810 ;
        RECT 67.560 76.910 68.460 77.810 ;
        RECT 62.960 76.010 67.860 76.310 ;
        RECT 113.670 75.860 119.270 76.260 ;
        RECT 124.070 75.560 124.870 76.960 ;
        RECT 120.170 74.660 124.870 75.560 ;
        RECT 127.070 76.260 127.970 77.160 ;
        RECT 133.470 76.260 134.370 77.160 ;
        RECT 128.870 75.360 133.770 75.660 ;
      LAYER met2 ;
        RECT 61.850 192.000 68.750 193.100 ;
        RECT 125.920 192.780 132.820 193.880 ;
        RECT 25.650 190.300 68.750 191.400 ;
        RECT 72.550 190.100 73.150 191.400 ;
        RECT 89.720 191.080 132.820 192.180 ;
        RECT 136.620 190.880 137.220 192.180 ;
        RECT 37.000 185.500 53.250 189.800 ;
        RECT 57.750 185.600 59.050 188.200 ;
        RECT 61.850 187.900 71.250 189.000 ;
        RECT 71.650 187.800 72.250 189.100 ;
        RECT 38.350 182.800 39.000 184.800 ;
        RECT 39.150 182.800 40.800 184.800 ;
        RECT 40.950 182.800 41.600 184.800 ;
        RECT 43.500 182.800 44.150 184.850 ;
        RECT 46.100 182.800 46.750 184.850 ;
        RECT 48.700 182.800 49.350 184.850 ;
        RECT 49.600 182.850 51.100 183.800 ;
        RECT 51.250 182.800 51.900 184.850 ;
        RECT 61.850 184.700 68.750 187.300 ;
        RECT 101.070 186.280 117.320 190.580 ;
        RECT 121.820 186.380 123.120 188.980 ;
        RECT 125.920 188.680 135.320 189.780 ;
        RECT 135.720 188.580 136.320 189.880 ;
        RECT 59.550 183.000 68.750 184.100 ;
        RECT 72.550 182.800 73.150 184.100 ;
        RECT 102.420 183.580 103.070 185.580 ;
        RECT 103.220 183.580 104.870 185.580 ;
        RECT 105.020 183.580 105.670 185.580 ;
        RECT 107.570 183.580 108.220 185.630 ;
        RECT 110.170 183.580 110.820 185.630 ;
        RECT 112.770 183.580 113.420 185.630 ;
        RECT 113.670 183.630 115.170 184.580 ;
        RECT 115.320 183.580 115.970 185.630 ;
        RECT 125.920 185.480 132.820 188.080 ;
        RECT 123.620 183.780 132.820 184.880 ;
        RECT 136.620 183.580 137.220 184.880 ;
        RECT 103.670 182.980 114.720 183.430 ;
        RECT 39.600 182.200 50.650 182.650 ;
        RECT 34.550 181.300 45.850 181.850 ;
        RECT 34.550 179.800 36.750 181.300 ;
        RECT 46.200 181.125 48.000 182.200 ;
        RECT 98.620 182.080 109.920 182.630 ;
        RECT 42.250 180.600 48.000 181.125 ;
        RECT 61.850 180.600 71.250 181.700 ;
        RECT 71.650 180.500 72.250 181.800 ;
        RECT 98.620 180.580 100.820 182.080 ;
        RECT 110.270 181.905 112.070 182.980 ;
        RECT 106.320 181.380 112.070 181.905 ;
        RECT 125.920 181.380 135.320 182.480 ;
        RECT 135.720 181.280 136.320 182.580 ;
        RECT 37.000 177.700 57.750 180.300 ;
        RECT 61.850 178.900 68.750 180.000 ;
        RECT 101.070 178.480 121.820 181.080 ;
        RECT 125.920 179.680 132.820 180.780 ;
        RECT 101.070 178.080 117.320 178.480 ;
        RECT 37.000 177.300 53.250 177.700 ;
        RECT 47.450 174.500 53.250 177.300 ;
        RECT 62.150 176.800 67.750 177.800 ;
        RECT 57.850 174.500 58.850 175.900 ;
        RECT 60.850 175.000 61.950 176.100 ;
        RECT 67.250 175.000 68.350 176.100 ;
        RECT 111.520 175.280 117.320 178.080 ;
        RECT 126.220 177.580 131.820 178.580 ;
        RECT 121.920 175.280 122.920 176.680 ;
        RECT 124.920 175.780 126.020 176.880 ;
        RECT 131.320 175.780 132.420 176.880 ;
        RECT 53.950 173.400 58.850 174.500 ;
        RECT 62.150 173.600 67.750 174.600 ;
        RECT 118.020 174.180 122.920 175.280 ;
        RECT 126.220 174.380 131.820 175.380 ;
        RECT 62.080 162.560 68.980 163.660 ;
        RECT 125.740 162.180 132.640 163.280 ;
        RECT 25.880 160.860 68.980 161.960 ;
        RECT 72.780 160.660 73.380 161.960 ;
        RECT 89.540 160.480 132.640 161.580 ;
        RECT 37.230 156.060 53.480 160.360 ;
        RECT 136.440 160.280 137.040 161.580 ;
        RECT 57.980 156.160 59.280 158.760 ;
        RECT 62.080 158.460 71.480 159.560 ;
        RECT 71.880 158.360 72.480 159.660 ;
        RECT 38.580 153.360 39.230 155.360 ;
        RECT 39.380 153.360 41.030 155.360 ;
        RECT 41.180 153.360 41.830 155.360 ;
        RECT 43.730 153.360 44.380 155.410 ;
        RECT 46.330 153.360 46.980 155.410 ;
        RECT 48.930 153.360 49.580 155.410 ;
        RECT 49.830 153.410 51.330 154.360 ;
        RECT 51.480 153.360 52.130 155.410 ;
        RECT 62.080 155.260 68.980 157.860 ;
        RECT 100.890 155.680 117.140 159.980 ;
        RECT 121.640 155.780 122.940 158.380 ;
        RECT 125.740 158.080 135.140 159.180 ;
        RECT 135.540 157.980 136.140 159.280 ;
        RECT 59.780 153.560 68.980 154.660 ;
        RECT 72.780 153.360 73.380 154.660 ;
        RECT 39.830 152.760 50.880 153.210 ;
        RECT 102.240 152.980 102.890 154.980 ;
        RECT 103.040 152.980 104.690 154.980 ;
        RECT 104.840 152.980 105.490 154.980 ;
        RECT 107.390 152.980 108.040 155.030 ;
        RECT 109.990 152.980 110.640 155.030 ;
        RECT 112.590 152.980 113.240 155.030 ;
        RECT 113.490 153.030 114.990 153.980 ;
        RECT 115.140 152.980 115.790 155.030 ;
        RECT 125.740 154.880 132.640 157.480 ;
        RECT 123.440 153.180 132.640 154.280 ;
        RECT 136.440 152.980 137.040 154.280 ;
        RECT 34.780 151.860 46.080 152.410 ;
        RECT 34.780 150.360 36.980 151.860 ;
        RECT 46.430 151.685 48.230 152.760 ;
        RECT 103.490 152.380 114.540 152.830 ;
        RECT 42.480 151.160 48.230 151.685 ;
        RECT 62.080 151.160 71.480 152.260 ;
        RECT 71.880 151.060 72.480 152.360 ;
        RECT 98.440 151.480 109.740 152.030 ;
        RECT 37.230 148.260 57.980 150.860 ;
        RECT 62.080 149.460 68.980 150.560 ;
        RECT 98.440 149.980 100.640 151.480 ;
        RECT 110.090 151.305 111.890 152.380 ;
        RECT 106.140 150.780 111.890 151.305 ;
        RECT 125.740 150.780 135.140 151.880 ;
        RECT 135.540 150.680 136.140 151.980 ;
        RECT 37.230 147.860 53.480 148.260 ;
        RECT 47.680 145.060 53.480 147.860 ;
        RECT 62.380 147.360 67.980 148.360 ;
        RECT 100.890 147.880 121.640 150.480 ;
        RECT 125.740 149.080 132.640 150.180 ;
        RECT 100.890 147.480 117.140 147.880 ;
        RECT 58.080 145.060 59.080 146.460 ;
        RECT 61.080 145.560 62.180 146.660 ;
        RECT 67.480 145.560 68.580 146.660 ;
        RECT 54.180 143.960 59.080 145.060 ;
        RECT 62.380 144.160 67.980 145.160 ;
        RECT 111.340 144.680 117.140 147.480 ;
        RECT 126.040 146.980 131.640 147.980 ;
        RECT 121.740 144.680 122.740 146.080 ;
        RECT 124.740 145.180 125.840 146.280 ;
        RECT 131.140 145.180 132.240 146.280 ;
        RECT 117.840 143.580 122.740 144.680 ;
        RECT 126.040 143.780 131.640 144.780 ;
        RECT 62.680 129.040 69.580 130.140 ;
        RECT 26.480 127.340 69.580 128.440 ;
        RECT 73.380 127.140 73.980 128.440 ;
        RECT 126.220 128.390 133.120 129.490 ;
        RECT 37.830 122.540 54.080 126.840 ;
        RECT 90.020 126.690 133.120 127.790 ;
        RECT 136.920 126.490 137.520 127.790 ;
        RECT 58.580 122.640 59.880 125.240 ;
        RECT 62.680 124.940 72.080 126.040 ;
        RECT 72.480 124.840 73.080 126.140 ;
        RECT 39.180 119.840 39.830 121.840 ;
        RECT 39.980 119.840 41.630 121.840 ;
        RECT 41.780 119.840 42.430 121.840 ;
        RECT 44.330 119.840 44.980 121.890 ;
        RECT 46.930 119.840 47.580 121.890 ;
        RECT 49.530 119.840 50.180 121.890 ;
        RECT 50.430 119.890 51.930 120.840 ;
        RECT 52.080 119.840 52.730 121.890 ;
        RECT 62.680 121.740 69.580 124.340 ;
        RECT 101.370 121.890 117.620 126.190 ;
        RECT 122.120 121.990 123.420 124.590 ;
        RECT 126.220 124.290 135.620 125.390 ;
        RECT 136.020 124.190 136.620 125.490 ;
        RECT 60.380 120.040 69.580 121.140 ;
        RECT 73.380 119.840 73.980 121.140 ;
        RECT 40.430 119.240 51.480 119.690 ;
        RECT 35.380 118.340 46.680 118.890 ;
        RECT 35.380 116.840 37.580 118.340 ;
        RECT 47.030 118.165 48.830 119.240 ;
        RECT 102.720 119.190 103.370 121.190 ;
        RECT 103.520 119.190 105.170 121.190 ;
        RECT 105.320 119.190 105.970 121.190 ;
        RECT 107.870 119.190 108.520 121.240 ;
        RECT 110.470 119.190 111.120 121.240 ;
        RECT 113.070 119.190 113.720 121.240 ;
        RECT 113.970 119.240 115.470 120.190 ;
        RECT 115.620 119.190 116.270 121.240 ;
        RECT 126.220 121.090 133.120 123.690 ;
        RECT 123.920 119.390 133.120 120.490 ;
        RECT 136.920 119.190 137.520 120.490 ;
        RECT 43.080 117.640 48.830 118.165 ;
        RECT 62.680 117.640 72.080 118.740 ;
        RECT 72.480 117.540 73.080 118.840 ;
        RECT 103.970 118.590 115.020 119.040 ;
        RECT 98.920 117.690 110.220 118.240 ;
        RECT 37.830 114.740 58.580 117.340 ;
        RECT 62.680 115.940 69.580 117.040 ;
        RECT 98.920 116.190 101.120 117.690 ;
        RECT 110.570 117.515 112.370 118.590 ;
        RECT 106.620 116.990 112.370 117.515 ;
        RECT 126.220 116.990 135.620 118.090 ;
        RECT 136.020 116.890 136.620 118.190 ;
        RECT 37.830 114.340 54.080 114.740 ;
        RECT 48.280 111.540 54.080 114.340 ;
        RECT 62.980 113.840 68.580 114.840 ;
        RECT 101.370 114.090 122.120 116.690 ;
        RECT 126.220 115.290 133.120 116.390 ;
        RECT 101.370 113.690 117.620 114.090 ;
        RECT 58.680 111.540 59.680 112.940 ;
        RECT 61.680 112.040 62.780 113.140 ;
        RECT 68.080 112.040 69.180 113.140 ;
        RECT 54.780 110.440 59.680 111.540 ;
        RECT 62.980 110.640 68.580 111.640 ;
        RECT 111.820 110.890 117.620 113.690 ;
        RECT 126.520 113.190 132.120 114.190 ;
        RECT 122.220 110.890 123.220 112.290 ;
        RECT 125.220 111.390 126.320 112.490 ;
        RECT 131.620 111.390 132.720 112.490 ;
        RECT 118.320 109.790 123.220 110.890 ;
        RECT 126.520 109.990 132.120 110.990 ;
        RECT 62.060 93.810 68.960 94.910 ;
        RECT 25.860 92.110 68.960 93.210 ;
        RECT 72.760 91.910 73.360 93.210 ;
        RECT 127.970 93.160 134.870 94.260 ;
        RECT 37.210 87.310 53.460 91.610 ;
        RECT 91.770 91.460 134.870 92.560 ;
        RECT 138.670 91.260 139.270 92.560 ;
        RECT 57.960 87.410 59.260 90.010 ;
        RECT 62.060 89.710 71.460 90.810 ;
        RECT 71.860 89.610 72.460 90.910 ;
        RECT 38.560 84.610 39.210 86.610 ;
        RECT 39.360 84.610 41.010 86.610 ;
        RECT 41.160 84.610 41.810 86.610 ;
        RECT 43.710 84.610 44.360 86.660 ;
        RECT 46.310 84.610 46.960 86.660 ;
        RECT 48.910 84.610 49.560 86.660 ;
        RECT 49.810 84.660 51.310 85.610 ;
        RECT 51.460 84.610 52.110 86.660 ;
        RECT 62.060 86.510 68.960 89.110 ;
        RECT 103.120 86.660 119.370 90.960 ;
        RECT 123.870 86.760 125.170 89.360 ;
        RECT 127.970 89.060 137.370 90.160 ;
        RECT 137.770 88.960 138.370 90.260 ;
        RECT 59.760 84.810 68.960 85.910 ;
        RECT 72.760 84.610 73.360 85.910 ;
        RECT 39.810 84.010 50.860 84.460 ;
        RECT 34.760 83.110 46.060 83.660 ;
        RECT 34.760 81.610 36.960 83.110 ;
        RECT 46.410 82.935 48.210 84.010 ;
        RECT 104.470 83.960 105.120 85.960 ;
        RECT 105.270 83.960 106.920 85.960 ;
        RECT 107.070 83.960 107.720 85.960 ;
        RECT 109.620 83.960 110.270 86.010 ;
        RECT 112.220 83.960 112.870 86.010 ;
        RECT 114.820 83.960 115.470 86.010 ;
        RECT 115.720 84.010 117.220 84.960 ;
        RECT 117.370 83.960 118.020 86.010 ;
        RECT 127.970 85.860 134.870 88.460 ;
        RECT 125.670 84.160 134.870 85.260 ;
        RECT 138.670 83.960 139.270 85.260 ;
        RECT 42.460 82.410 48.210 82.935 ;
        RECT 62.060 82.410 71.460 83.510 ;
        RECT 71.860 82.310 72.460 83.610 ;
        RECT 105.720 83.360 116.770 83.810 ;
        RECT 100.670 82.460 111.970 83.010 ;
        RECT 37.210 79.510 57.960 82.110 ;
        RECT 62.060 80.710 68.960 81.810 ;
        RECT 100.670 80.960 102.870 82.460 ;
        RECT 112.320 82.285 114.120 83.360 ;
        RECT 108.370 81.760 114.120 82.285 ;
        RECT 127.970 81.760 137.370 82.860 ;
        RECT 137.770 81.660 138.370 82.960 ;
        RECT 37.210 79.110 53.460 79.510 ;
        RECT 47.660 76.310 53.460 79.110 ;
        RECT 62.360 78.610 67.960 79.610 ;
        RECT 103.120 78.860 123.870 81.460 ;
        RECT 127.970 80.060 134.870 81.160 ;
        RECT 103.120 78.460 119.370 78.860 ;
        RECT 58.060 76.310 59.060 77.710 ;
        RECT 61.060 76.810 62.160 77.910 ;
        RECT 67.460 76.810 68.560 77.910 ;
        RECT 54.160 75.210 59.060 76.310 ;
        RECT 62.360 75.410 67.960 76.410 ;
        RECT 113.570 75.660 119.370 78.460 ;
        RECT 128.270 77.960 133.870 78.960 ;
        RECT 123.970 75.660 124.970 77.060 ;
        RECT 126.970 76.160 128.070 77.260 ;
        RECT 133.370 76.160 134.470 77.260 ;
        RECT 120.070 74.560 124.970 75.660 ;
        RECT 128.270 74.760 133.870 75.760 ;
      LAYER via2 ;
        RECT 62.550 192.100 64.150 193.000 ;
        RECT 126.620 192.880 128.220 193.780 ;
        RECT 25.750 190.400 27.250 191.300 ;
        RECT 72.650 190.200 73.050 191.300 ;
        RECT 89.820 191.180 91.320 192.080 ;
        RECT 136.720 190.980 137.120 192.080 ;
        RECT 37.050 185.550 53.200 186.900 ;
        RECT 57.850 185.700 58.950 188.100 ;
        RECT 69.750 188.000 71.150 188.900 ;
        RECT 71.750 187.900 72.150 189.000 ;
        RECT 38.400 182.850 38.950 183.200 ;
        RECT 39.200 183.650 40.550 184.750 ;
        RECT 41.000 184.400 41.550 184.750 ;
        RECT 43.550 182.850 44.100 183.200 ;
        RECT 46.150 184.400 46.700 184.750 ;
        RECT 51.300 184.400 51.850 184.750 ;
        RECT 67.350 184.800 68.250 187.200 ;
        RECT 101.120 186.330 117.270 187.680 ;
        RECT 121.920 186.480 123.020 188.880 ;
        RECT 133.820 188.780 135.220 189.680 ;
        RECT 135.820 188.680 136.220 189.780 ;
        RECT 48.750 182.850 49.300 183.200 ;
        RECT 49.700 182.900 51.050 183.750 ;
        RECT 59.650 183.100 60.650 184.000 ;
        RECT 72.650 182.900 73.050 184.000 ;
        RECT 102.470 183.630 103.020 183.980 ;
        RECT 103.270 184.430 104.620 185.530 ;
        RECT 105.070 185.180 105.620 185.530 ;
        RECT 107.620 183.630 108.170 183.980 ;
        RECT 110.220 185.180 110.770 185.530 ;
        RECT 115.370 185.180 115.920 185.530 ;
        RECT 131.420 185.580 132.320 187.980 ;
        RECT 112.820 183.630 113.370 183.980 ;
        RECT 113.770 183.680 115.120 184.530 ;
        RECT 123.720 183.880 124.720 184.780 ;
        RECT 136.720 183.680 137.120 184.780 ;
        RECT 69.750 180.700 71.150 181.600 ;
        RECT 71.750 180.600 72.150 181.700 ;
        RECT 133.820 181.480 135.220 182.380 ;
        RECT 135.820 181.380 136.220 182.480 ;
        RECT 37.100 179.050 53.150 180.300 ;
        RECT 62.150 179.000 64.150 179.900 ;
        RECT 101.170 179.830 117.220 181.080 ;
        RECT 126.220 179.780 128.220 180.680 ;
        RECT 64.750 176.900 66.650 177.700 ;
        RECT 57.950 174.400 58.750 175.800 ;
        RECT 54.050 173.500 58.750 174.400 ;
        RECT 60.950 175.100 61.850 176.000 ;
        RECT 67.350 175.100 68.250 176.000 ;
        RECT 128.820 177.680 130.720 178.480 ;
        RECT 122.020 175.180 122.820 176.580 ;
        RECT 62.550 173.700 64.150 174.500 ;
        RECT 118.120 174.280 122.820 175.180 ;
        RECT 125.020 175.880 125.920 176.780 ;
        RECT 131.420 175.880 132.320 176.780 ;
        RECT 126.620 174.480 128.220 175.280 ;
        RECT 62.780 162.660 64.380 163.560 ;
        RECT 126.440 162.280 128.040 163.180 ;
        RECT 25.980 160.960 27.480 161.860 ;
        RECT 72.880 160.760 73.280 161.860 ;
        RECT 89.640 160.580 91.140 161.480 ;
        RECT 136.540 160.380 136.940 161.480 ;
        RECT 37.280 156.110 53.430 157.460 ;
        RECT 58.080 156.260 59.180 158.660 ;
        RECT 69.980 158.560 71.380 159.460 ;
        RECT 71.980 158.460 72.380 159.560 ;
        RECT 38.630 153.410 39.180 153.760 ;
        RECT 39.430 154.210 40.780 155.310 ;
        RECT 41.230 154.960 41.780 155.310 ;
        RECT 43.780 153.410 44.330 153.760 ;
        RECT 46.380 154.960 46.930 155.310 ;
        RECT 51.530 154.960 52.080 155.310 ;
        RECT 67.580 155.360 68.480 157.760 ;
        RECT 100.940 155.730 117.090 157.080 ;
        RECT 121.740 155.880 122.840 158.280 ;
        RECT 133.640 158.180 135.040 159.080 ;
        RECT 135.640 158.080 136.040 159.180 ;
        RECT 48.980 153.410 49.530 153.760 ;
        RECT 49.930 153.460 51.280 154.310 ;
        RECT 59.880 153.660 60.880 154.560 ;
        RECT 72.880 153.460 73.280 154.560 ;
        RECT 102.290 153.030 102.840 153.380 ;
        RECT 103.090 153.830 104.440 154.930 ;
        RECT 104.890 154.580 105.440 154.930 ;
        RECT 107.440 153.030 107.990 153.380 ;
        RECT 110.040 154.580 110.590 154.930 ;
        RECT 115.190 154.580 115.740 154.930 ;
        RECT 131.240 154.980 132.140 157.380 ;
        RECT 112.640 153.030 113.190 153.380 ;
        RECT 113.590 153.080 114.940 153.930 ;
        RECT 123.540 153.280 124.540 154.180 ;
        RECT 136.540 153.080 136.940 154.180 ;
        RECT 69.980 151.260 71.380 152.160 ;
        RECT 71.980 151.160 72.380 152.260 ;
        RECT 37.330 149.610 53.380 150.860 ;
        RECT 62.380 149.560 64.380 150.460 ;
        RECT 133.640 150.880 135.040 151.780 ;
        RECT 135.640 150.780 136.040 151.880 ;
        RECT 100.990 149.230 117.040 150.480 ;
        RECT 64.980 147.460 66.880 148.260 ;
        RECT 126.040 149.180 128.040 150.080 ;
        RECT 58.180 144.960 58.980 146.360 ;
        RECT 54.280 144.060 58.980 144.960 ;
        RECT 61.180 145.660 62.080 146.560 ;
        RECT 67.580 145.660 68.480 146.560 ;
        RECT 62.780 144.260 64.380 145.060 ;
        RECT 128.640 147.080 130.540 147.880 ;
        RECT 121.840 144.580 122.640 145.980 ;
        RECT 117.940 143.680 122.640 144.580 ;
        RECT 124.840 145.280 125.740 146.180 ;
        RECT 131.240 145.280 132.140 146.180 ;
        RECT 126.440 143.880 128.040 144.680 ;
        RECT 63.380 129.140 64.980 130.040 ;
        RECT 126.920 128.490 128.520 129.390 ;
        RECT 26.580 127.440 28.080 128.340 ;
        RECT 73.480 127.240 73.880 128.340 ;
        RECT 90.120 126.790 91.620 127.690 ;
        RECT 137.020 126.590 137.420 127.690 ;
        RECT 37.880 122.590 54.030 123.940 ;
        RECT 58.680 122.740 59.780 125.140 ;
        RECT 70.580 125.040 71.980 125.940 ;
        RECT 72.580 124.940 72.980 126.040 ;
        RECT 39.230 119.890 39.780 120.240 ;
        RECT 40.030 120.690 41.380 121.790 ;
        RECT 41.830 121.440 42.380 121.790 ;
        RECT 44.380 119.890 44.930 120.240 ;
        RECT 46.980 121.440 47.530 121.790 ;
        RECT 52.130 121.440 52.680 121.790 ;
        RECT 68.180 121.840 69.080 124.240 ;
        RECT 101.420 121.940 117.570 123.290 ;
        RECT 122.220 122.090 123.320 124.490 ;
        RECT 134.120 124.390 135.520 125.290 ;
        RECT 136.120 124.290 136.520 125.390 ;
        RECT 49.580 119.890 50.130 120.240 ;
        RECT 50.530 119.940 51.880 120.790 ;
        RECT 60.480 120.140 61.480 121.040 ;
        RECT 73.480 119.940 73.880 121.040 ;
        RECT 102.770 119.240 103.320 119.590 ;
        RECT 103.570 120.040 104.920 121.140 ;
        RECT 105.370 120.790 105.920 121.140 ;
        RECT 107.920 119.240 108.470 119.590 ;
        RECT 110.520 120.790 111.070 121.140 ;
        RECT 115.670 120.790 116.220 121.140 ;
        RECT 131.720 121.190 132.620 123.590 ;
        RECT 113.120 119.240 113.670 119.590 ;
        RECT 114.070 119.290 115.420 120.140 ;
        RECT 124.020 119.490 125.020 120.390 ;
        RECT 137.020 119.290 137.420 120.390 ;
        RECT 70.580 117.740 71.980 118.640 ;
        RECT 72.580 117.640 72.980 118.740 ;
        RECT 37.930 116.090 53.980 117.340 ;
        RECT 62.980 116.040 64.980 116.940 ;
        RECT 134.120 117.090 135.520 117.990 ;
        RECT 136.120 116.990 136.520 118.090 ;
        RECT 101.470 115.440 117.520 116.690 ;
        RECT 65.580 113.940 67.480 114.740 ;
        RECT 126.520 115.390 128.520 116.290 ;
        RECT 58.780 111.440 59.580 112.840 ;
        RECT 54.880 110.540 59.580 111.440 ;
        RECT 61.780 112.140 62.680 113.040 ;
        RECT 68.180 112.140 69.080 113.040 ;
        RECT 63.380 110.740 64.980 111.540 ;
        RECT 129.120 113.290 131.020 114.090 ;
        RECT 122.320 110.790 123.120 112.190 ;
        RECT 118.420 109.890 123.120 110.790 ;
        RECT 125.320 111.490 126.220 112.390 ;
        RECT 131.720 111.490 132.620 112.390 ;
        RECT 126.920 110.090 128.520 110.890 ;
        RECT 62.760 93.910 64.360 94.810 ;
        RECT 128.670 93.260 130.270 94.160 ;
        RECT 25.960 92.210 27.460 93.110 ;
        RECT 72.860 92.010 73.260 93.110 ;
        RECT 91.870 91.560 93.370 92.460 ;
        RECT 138.770 91.360 139.170 92.460 ;
        RECT 37.260 87.360 53.410 88.710 ;
        RECT 58.060 87.510 59.160 89.910 ;
        RECT 69.960 89.810 71.360 90.710 ;
        RECT 71.960 89.710 72.360 90.810 ;
        RECT 38.610 84.660 39.160 85.010 ;
        RECT 39.410 85.460 40.760 86.560 ;
        RECT 41.210 86.210 41.760 86.560 ;
        RECT 43.760 84.660 44.310 85.010 ;
        RECT 46.360 86.210 46.910 86.560 ;
        RECT 51.510 86.210 52.060 86.560 ;
        RECT 67.560 86.610 68.460 89.010 ;
        RECT 103.170 86.710 119.320 88.060 ;
        RECT 123.970 86.860 125.070 89.260 ;
        RECT 135.870 89.160 137.270 90.060 ;
        RECT 137.870 89.060 138.270 90.160 ;
        RECT 48.960 84.660 49.510 85.010 ;
        RECT 49.910 84.710 51.260 85.560 ;
        RECT 59.860 84.910 60.860 85.810 ;
        RECT 72.860 84.710 73.260 85.810 ;
        RECT 104.520 84.010 105.070 84.360 ;
        RECT 105.320 84.810 106.670 85.910 ;
        RECT 107.120 85.560 107.670 85.910 ;
        RECT 109.670 84.010 110.220 84.360 ;
        RECT 112.270 85.560 112.820 85.910 ;
        RECT 117.420 85.560 117.970 85.910 ;
        RECT 133.470 85.960 134.370 88.360 ;
        RECT 114.870 84.010 115.420 84.360 ;
        RECT 115.820 84.060 117.170 84.910 ;
        RECT 125.770 84.260 126.770 85.160 ;
        RECT 138.770 84.060 139.170 85.160 ;
        RECT 69.960 82.510 71.360 83.410 ;
        RECT 71.960 82.410 72.360 83.510 ;
        RECT 37.310 80.860 53.360 82.110 ;
        RECT 62.360 80.810 64.360 81.710 ;
        RECT 135.870 81.860 137.270 82.760 ;
        RECT 137.870 81.760 138.270 82.860 ;
        RECT 103.220 80.210 119.270 81.460 ;
        RECT 64.960 78.710 66.860 79.510 ;
        RECT 128.270 80.160 130.270 81.060 ;
        RECT 58.160 76.210 58.960 77.610 ;
        RECT 54.260 75.310 58.960 76.210 ;
        RECT 61.160 76.910 62.060 77.810 ;
        RECT 67.560 76.910 68.460 77.810 ;
        RECT 62.760 75.510 64.360 76.310 ;
        RECT 130.870 78.060 132.770 78.860 ;
        RECT 124.070 75.560 124.870 76.960 ;
        RECT 120.170 74.660 124.870 75.560 ;
        RECT 127.070 76.260 127.970 77.160 ;
        RECT 133.470 76.260 134.370 77.160 ;
        RECT 128.670 74.860 130.270 75.660 ;
      LAYER met3 ;
        RECT 57.410 222.475 150.750 222.940 ;
        RECT 148.400 222.470 150.750 222.475 ;
        RECT 60.255 221.460 150.700 221.930 ;
        RECT 63.025 220.440 150.810 220.910 ;
        RECT 58.795 219.310 150.700 219.780 ;
        RECT 61.705 218.170 150.750 218.640 ;
        RECT 61.855 217.150 150.640 217.620 ;
        RECT 57.695 216.230 150.700 216.700 ;
        RECT 60.255 215.370 150.590 215.840 ;
        RECT 89.720 195.600 91.420 195.680 ;
        RECT 12.450 194.900 27.310 195.060 ;
        RECT 12.450 192.980 27.350 194.900 ;
        RECT 12.450 11.980 14.530 192.980 ;
        RECT 25.650 185.100 27.350 192.980 ;
        RECT 27.950 185.500 56.450 189.800 ;
        RECT 57.750 185.400 59.050 188.200 ;
        RECT 25.650 183.600 40.600 185.100 ;
        RECT 57.750 184.900 60.750 185.400 ;
        RECT 50.050 184.800 60.750 184.900 ;
        RECT 37.250 183.550 40.600 183.600 ;
        RECT 40.900 184.400 60.750 184.800 ;
        RECT 40.900 184.350 51.900 184.400 ;
        RECT 40.900 183.550 49.200 184.350 ;
        RECT 49.650 184.000 53.000 184.050 ;
        RECT 38.350 182.800 49.350 183.250 ;
        RECT 41.050 182.000 49.350 182.800 ;
        RECT 49.650 182.100 58.850 184.000 ;
        RECT 59.550 183.000 60.750 184.400 ;
        RECT 27.950 175.800 56.450 180.450 ;
        RECT 57.850 174.500 58.850 182.100 ;
        RECT 62.450 180.200 64.250 195.600 ;
        RECT 69.650 194.000 91.420 195.600 ;
        RECT 60.850 178.600 64.250 180.200 ;
        RECT 60.850 175.000 61.950 178.600 ;
        RECT 53.950 173.400 58.850 174.500 ;
        RECT 62.450 173.600 64.250 177.800 ;
        RECT 64.650 176.800 66.750 189.800 ;
        RECT 67.250 175.000 68.350 187.300 ;
        RECT 69.650 180.600 71.250 194.000 ;
        RECT 71.650 175.800 72.250 189.100 ;
        RECT 72.550 182.800 73.150 191.400 ;
        RECT 89.720 185.880 91.420 194.000 ;
        RECT 92.020 186.280 120.520 190.580 ;
        RECT 121.820 186.180 123.120 188.980 ;
        RECT 89.720 184.380 104.670 185.880 ;
        RECT 121.820 185.680 124.820 186.180 ;
        RECT 114.120 185.580 124.820 185.680 ;
        RECT 101.320 184.330 104.670 184.380 ;
        RECT 104.970 185.180 124.820 185.580 ;
        RECT 104.970 185.130 115.970 185.180 ;
        RECT 104.970 184.330 113.270 185.130 ;
        RECT 113.720 184.780 117.070 184.830 ;
        RECT 102.420 183.580 113.420 184.030 ;
        RECT 105.120 182.780 113.420 183.580 ;
        RECT 113.720 182.880 122.920 184.780 ;
        RECT 123.620 183.780 124.820 185.180 ;
        RECT 92.020 176.580 120.520 181.230 ;
        RECT 121.920 175.280 122.920 182.880 ;
        RECT 126.520 180.980 128.320 196.380 ;
        RECT 133.720 196.345 135.320 196.380 ;
        RECT 146.675 196.345 148.290 196.360 ;
        RECT 133.720 194.755 148.290 196.345 ;
        RECT 124.920 179.380 128.320 180.980 ;
        RECT 124.920 175.780 126.020 179.380 ;
        RECT 118.020 174.180 122.920 175.280 ;
        RECT 126.520 174.380 128.320 178.580 ;
        RECT 128.720 177.580 130.820 190.580 ;
        RECT 131.320 175.780 132.420 188.080 ;
        RECT 133.720 181.380 135.320 194.755 ;
        RECT 135.720 176.580 136.320 189.880 ;
        RECT 136.620 183.580 137.220 192.180 ;
        RECT 146.675 172.590 148.290 194.755 ;
        RECT 25.450 170.990 148.290 172.590 ;
        RECT 25.460 163.340 27.595 170.990 ;
        RECT 146.675 170.985 148.290 170.990 ;
        RECT 25.470 161.840 27.580 163.340 ;
        RECT 25.880 155.660 27.580 161.840 ;
        RECT 28.180 156.060 56.680 160.360 ;
        RECT 57.980 155.960 59.280 158.760 ;
        RECT 25.880 154.160 40.830 155.660 ;
        RECT 57.980 155.460 60.980 155.960 ;
        RECT 50.280 155.360 60.980 155.460 ;
        RECT 37.480 154.110 40.830 154.160 ;
        RECT 41.130 154.960 60.980 155.360 ;
        RECT 41.130 154.910 52.130 154.960 ;
        RECT 41.130 154.110 49.430 154.910 ;
        RECT 49.880 154.560 53.230 154.610 ;
        RECT 38.580 153.360 49.580 153.810 ;
        RECT 41.280 152.560 49.580 153.360 ;
        RECT 49.880 152.660 59.080 154.560 ;
        RECT 59.780 153.560 60.980 154.960 ;
        RECT 28.180 146.360 56.680 151.010 ;
        RECT 58.080 145.060 59.080 152.660 ;
        RECT 62.680 150.760 64.480 166.160 ;
        RECT 69.880 164.970 71.480 166.160 ;
        RECT 89.540 164.970 91.240 165.080 ;
        RECT 69.880 163.270 91.240 164.970 ;
        RECT 61.080 149.160 64.480 150.760 ;
        RECT 61.080 145.560 62.180 149.160 ;
        RECT 54.180 143.960 59.080 145.060 ;
        RECT 62.680 144.160 64.480 148.360 ;
        RECT 64.880 147.360 66.980 160.360 ;
        RECT 67.480 145.560 68.580 157.860 ;
        RECT 69.880 151.160 71.480 163.270 ;
        RECT 71.880 146.360 72.480 159.660 ;
        RECT 72.780 153.360 73.380 161.960 ;
        RECT 89.540 155.280 91.240 163.270 ;
        RECT 91.840 155.680 120.340 159.980 ;
        RECT 121.640 155.580 122.940 158.380 ;
        RECT 89.540 153.780 104.490 155.280 ;
        RECT 121.640 155.080 124.640 155.580 ;
        RECT 113.940 154.980 124.640 155.080 ;
        RECT 101.140 153.730 104.490 153.780 ;
        RECT 104.790 154.580 124.640 154.980 ;
        RECT 104.790 154.530 115.790 154.580 ;
        RECT 104.790 153.730 113.090 154.530 ;
        RECT 113.540 154.180 116.890 154.230 ;
        RECT 102.240 152.980 113.240 153.430 ;
        RECT 104.940 152.180 113.240 152.980 ;
        RECT 113.540 152.280 122.740 154.180 ;
        RECT 123.440 153.180 124.640 154.580 ;
        RECT 91.840 145.980 120.340 150.630 ;
        RECT 121.740 144.680 122.740 152.280 ;
        RECT 126.340 150.380 128.140 165.780 ;
        RECT 133.540 164.180 147.610 165.780 ;
        RECT 124.740 148.780 128.140 150.380 ;
        RECT 124.740 145.180 125.840 148.780 ;
        RECT 117.840 143.580 122.740 144.680 ;
        RECT 126.340 143.780 128.140 147.980 ;
        RECT 128.540 146.980 130.640 159.980 ;
        RECT 131.140 145.180 132.240 157.480 ;
        RECT 133.540 150.780 135.140 164.180 ;
        RECT 135.540 145.980 136.140 159.280 ;
        RECT 136.440 152.980 137.040 161.580 ;
        RECT 146.020 141.990 147.600 164.180 ;
        RECT 26.450 140.410 147.600 141.990 ;
        RECT 26.480 122.140 28.180 140.410 ;
        RECT 28.780 122.540 57.280 126.840 ;
        RECT 58.580 122.440 59.880 125.240 ;
        RECT 26.480 120.640 41.430 122.140 ;
        RECT 58.580 121.940 61.580 122.440 ;
        RECT 50.880 121.840 61.580 121.940 ;
        RECT 38.080 120.590 41.430 120.640 ;
        RECT 41.730 121.440 61.580 121.840 ;
        RECT 41.730 121.390 52.730 121.440 ;
        RECT 41.730 120.590 50.030 121.390 ;
        RECT 50.480 121.040 53.830 121.090 ;
        RECT 39.180 119.840 50.180 120.290 ;
        RECT 41.880 119.040 50.180 119.840 ;
        RECT 50.480 119.140 59.680 121.040 ;
        RECT 60.380 120.040 61.580 121.440 ;
        RECT 28.780 112.840 57.280 117.490 ;
        RECT 58.680 111.540 59.680 119.140 ;
        RECT 63.280 117.240 65.080 132.640 ;
        RECT 70.480 131.400 72.080 132.640 ;
        RECT 70.480 129.800 91.830 131.400 ;
        RECT 61.680 115.640 65.080 117.240 ;
        RECT 61.680 112.040 62.780 115.640 ;
        RECT 54.780 110.440 59.680 111.540 ;
        RECT 63.280 110.640 65.080 114.840 ;
        RECT 65.480 113.840 67.580 126.840 ;
        RECT 68.080 112.040 69.180 124.340 ;
        RECT 70.480 117.640 72.080 129.800 ;
        RECT 72.480 112.840 73.080 126.140 ;
        RECT 73.380 119.840 73.980 128.440 ;
        RECT 90.020 121.490 91.720 129.800 ;
        RECT 92.320 121.890 120.820 126.190 ;
        RECT 122.120 121.790 123.420 124.590 ;
        RECT 90.020 119.990 104.970 121.490 ;
        RECT 122.120 121.290 125.120 121.790 ;
        RECT 114.420 121.190 125.120 121.290 ;
        RECT 101.620 119.940 104.970 119.990 ;
        RECT 105.270 120.790 125.120 121.190 ;
        RECT 105.270 120.740 116.270 120.790 ;
        RECT 105.270 119.940 113.570 120.740 ;
        RECT 114.020 120.390 117.370 120.440 ;
        RECT 102.720 119.190 113.720 119.640 ;
        RECT 105.420 118.390 113.720 119.190 ;
        RECT 114.020 118.490 123.220 120.390 ;
        RECT 123.920 119.390 125.120 120.790 ;
        RECT 92.320 112.190 120.820 116.840 ;
        RECT 122.220 110.890 123.220 118.490 ;
        RECT 126.820 116.590 128.620 131.990 ;
        RECT 134.020 131.330 135.620 131.990 ;
        RECT 134.020 129.730 146.800 131.330 ;
        RECT 125.220 114.990 128.620 116.590 ;
        RECT 125.220 111.390 126.320 114.990 ;
        RECT 118.320 109.790 123.220 110.890 ;
        RECT 126.820 109.990 128.620 114.190 ;
        RECT 129.020 113.190 131.120 126.190 ;
        RECT 131.620 111.390 132.720 123.690 ;
        RECT 134.020 116.990 135.620 129.730 ;
        RECT 136.020 112.190 136.620 125.490 ;
        RECT 136.920 119.190 137.520 127.790 ;
        RECT 25.860 108.370 27.560 108.450 ;
        RECT 145.200 108.370 146.800 129.730 ;
        RECT 25.860 106.770 146.800 108.370 ;
        RECT 25.860 86.910 27.560 106.770 ;
        RECT 28.160 87.310 56.660 91.610 ;
        RECT 57.960 87.210 59.260 90.010 ;
        RECT 25.860 85.410 40.810 86.910 ;
        RECT 57.960 86.710 60.960 87.210 ;
        RECT 50.260 86.610 60.960 86.710 ;
        RECT 37.460 85.360 40.810 85.410 ;
        RECT 41.110 86.210 60.960 86.610 ;
        RECT 41.110 86.160 52.110 86.210 ;
        RECT 41.110 85.360 49.410 86.160 ;
        RECT 49.860 85.810 53.210 85.860 ;
        RECT 38.560 84.610 49.560 85.060 ;
        RECT 41.260 83.810 49.560 84.610 ;
        RECT 49.860 83.910 59.060 85.810 ;
        RECT 59.760 84.810 60.960 86.210 ;
        RECT 28.160 77.610 56.660 82.260 ;
        RECT 58.060 76.310 59.060 83.910 ;
        RECT 62.660 82.010 64.460 97.410 ;
        RECT 69.860 97.280 71.460 97.410 ;
        RECT 69.860 96.060 93.440 97.280 ;
        RECT 69.860 95.680 93.470 96.060 ;
        RECT 61.060 80.410 64.460 82.010 ;
        RECT 61.060 76.810 62.160 80.410 ;
        RECT 54.160 75.210 59.060 76.310 ;
        RECT 62.660 75.410 64.460 79.610 ;
        RECT 64.860 78.610 66.960 91.610 ;
        RECT 67.460 76.810 68.560 89.110 ;
        RECT 69.860 82.410 71.460 95.680 ;
        RECT 71.860 77.610 72.460 90.910 ;
        RECT 72.760 84.610 73.360 93.210 ;
        RECT 91.770 86.260 93.470 95.680 ;
        RECT 94.070 86.660 122.570 90.960 ;
        RECT 123.870 86.560 125.170 89.360 ;
        RECT 91.770 84.760 106.720 86.260 ;
        RECT 123.870 86.060 126.870 86.560 ;
        RECT 116.170 85.960 126.870 86.060 ;
        RECT 103.370 84.710 106.720 84.760 ;
        RECT 107.020 85.560 126.870 85.960 ;
        RECT 107.020 85.510 118.020 85.560 ;
        RECT 107.020 84.710 115.320 85.510 ;
        RECT 115.770 85.160 119.120 85.210 ;
        RECT 104.470 83.960 115.470 84.410 ;
        RECT 107.170 83.160 115.470 83.960 ;
        RECT 115.770 83.260 124.970 85.160 ;
        RECT 125.670 84.160 126.870 85.560 ;
        RECT 94.070 76.960 122.570 81.610 ;
        RECT 123.970 75.660 124.970 83.260 ;
        RECT 128.570 81.360 130.370 96.760 ;
        RECT 135.770 95.160 148.200 96.760 ;
        RECT 126.970 79.760 130.370 81.360 ;
        RECT 126.970 76.160 128.070 79.760 ;
        RECT 120.070 74.560 124.970 75.660 ;
        RECT 128.570 74.760 130.370 78.960 ;
        RECT 130.770 77.960 132.870 90.960 ;
        RECT 133.370 76.160 134.470 88.460 ;
        RECT 135.770 81.760 137.370 95.160 ;
        RECT 137.770 76.960 138.370 90.260 ;
        RECT 138.670 83.960 139.270 92.560 ;
        RECT 146.625 7.210 148.180 95.160 ;
        RECT 134.380 5.655 148.180 7.210 ;
      LAYER via3 ;
        RECT 28.250 185.800 56.050 189.500 ;
        RECT 28.250 176.100 56.150 180.200 ;
        RECT 64.750 185.600 66.650 189.700 ;
        RECT 62.550 175.900 64.150 177.700 ;
        RECT 72.650 185.600 73.050 189.700 ;
        RECT 92.320 186.580 120.120 190.280 ;
        RECT 71.750 175.900 72.150 180.400 ;
        RECT 92.320 176.880 120.220 180.980 ;
        RECT 128.820 186.380 130.720 190.480 ;
        RECT 126.620 176.680 128.220 178.480 ;
        RECT 136.720 186.380 137.120 190.480 ;
        RECT 135.820 176.680 136.220 181.180 ;
        RECT 28.480 156.360 56.280 160.060 ;
        RECT 28.480 146.660 56.380 150.760 ;
        RECT 64.980 156.160 66.880 160.260 ;
        RECT 62.780 146.460 64.380 148.260 ;
        RECT 72.880 156.160 73.280 160.260 ;
        RECT 92.140 155.980 119.940 159.680 ;
        RECT 71.980 146.460 72.380 150.960 ;
        RECT 92.140 146.280 120.040 150.380 ;
        RECT 128.640 155.780 130.540 159.880 ;
        RECT 126.440 146.080 128.040 147.880 ;
        RECT 136.540 155.780 136.940 159.880 ;
        RECT 135.640 146.080 136.040 150.580 ;
        RECT 29.080 122.840 56.880 126.540 ;
        RECT 29.080 113.140 56.980 117.240 ;
        RECT 65.580 122.640 67.480 126.740 ;
        RECT 63.380 112.940 64.980 114.740 ;
        RECT 73.480 122.640 73.880 126.740 ;
        RECT 92.620 122.190 120.420 125.890 ;
        RECT 72.580 112.940 72.980 117.440 ;
        RECT 92.620 112.490 120.520 116.590 ;
        RECT 129.120 121.990 131.020 126.090 ;
        RECT 126.920 112.290 128.520 114.090 ;
        RECT 137.020 121.990 137.420 126.090 ;
        RECT 136.120 112.290 136.520 116.790 ;
        RECT 28.460 87.610 56.260 91.310 ;
        RECT 28.460 77.910 56.360 82.010 ;
        RECT 64.960 87.410 66.860 91.510 ;
        RECT 62.760 77.710 64.360 79.510 ;
        RECT 72.860 87.410 73.260 91.510 ;
        RECT 94.370 86.960 122.170 90.660 ;
        RECT 71.960 77.710 72.360 82.210 ;
        RECT 94.370 77.260 122.270 81.360 ;
        RECT 130.870 86.760 132.770 90.860 ;
        RECT 128.670 77.060 130.270 78.860 ;
        RECT 138.770 86.760 139.170 90.860 ;
        RECT 137.870 77.060 138.270 81.560 ;
        RECT 12.530 12.500 14.440 13.000 ;
        RECT 134.550 5.730 135.010 7.150 ;
      LAYER met4 ;
        RECT 121.750 214.950 122.050 224.760 ;
        RECT 125.430 214.910 125.730 224.760 ;
        RECT 129.110 215.070 129.410 224.760 ;
        RECT 132.790 215.120 133.090 224.760 ;
        RECT 136.470 214.610 136.770 224.760 ;
        RECT 140.150 214.860 140.450 224.760 ;
        RECT 143.830 215.120 144.130 224.760 ;
        RECT 147.510 214.960 147.810 224.760 ;
        RECT 6.500 185.000 144.000 193.000 ;
        RECT 27.000 175.000 157.530 182.000 ;
        RECT 6.500 155.000 144.000 163.000 ;
        RECT 27.000 145.000 157.530 152.000 ;
        RECT 6.500 120.000 144.000 128.000 ;
        RECT 27.000 111.000 157.530 118.000 ;
        RECT 6.500 86.000 144.000 92.000 ;
        RECT 27.000 77.000 157.530 84.000 ;
        RECT 94.070 76.960 141.970 77.000 ;
        RECT 12.085 12.455 142.625 13.045 ;
        RECT 134.480 1.000 135.080 7.280 ;
        RECT 142.035 2.410 142.625 12.455 ;
        RECT 142.030 1.810 157.160 2.410 ;
        RECT 156.560 1.000 157.160 1.810 ;
  END
END tt_um_guitar_pedal
END LIBRARY

