** sch_path: /home/ttuser/pdk/sky130A/libs.tech/xschem/tgate.sch
**.subckt tgate IN OUT CTRL CTRLB
*.ipin IN
*.opin OUT
*.ipin CTRL
*.ipin CTRLB
XM11 OUT CTRLB IN IN sky130_fd_pr__pfet_01v8 L=1 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 IN CTRL OUT OUT sky130_fd_pr__nfet_01v8 L=1 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
**.ends
.end
