magic
tech sky130A
magscale 1 2
timestamp 1713492510
<< metal2 >>
rect 14960 44600 15140 44620
rect 14960 44480 14980 44600
rect 15120 44480 15140 44600
rect 14960 44460 15140 44480
rect 15000 39944 15100 44460
rect 17380 44400 17600 44420
rect 17380 44280 17400 44400
rect 17580 44280 17600 44400
rect 17380 44260 17600 44280
rect 15380 44200 15600 44220
rect 15380 44040 15400 44200
rect 15580 44040 15600 44200
rect 15380 44020 15600 44040
rect 12644 39844 15100 39944
rect 12644 39108 12744 39844
rect 12644 38710 12656 39108
rect 12734 38710 12744 39108
rect 12644 38698 12744 38710
rect 15440 33936 15540 44020
rect 17080 44000 17320 44020
rect 17080 43820 17100 44000
rect 17300 43820 17320 44000
rect 17080 43800 17320 43820
rect 15760 43780 15980 43800
rect 15760 43620 15780 43780
rect 15960 43620 15980 43780
rect 15760 43600 15980 43620
rect 15820 38120 15920 43600
rect 16820 43540 17000 43560
rect 16820 43420 16840 43540
rect 16980 43420 17000 43540
rect 16820 43400 17000 43420
rect 16080 43340 16260 43360
rect 16080 43220 16100 43340
rect 16240 43220 16260 43340
rect 16080 43200 16260 43220
rect 12694 33836 15540 33936
rect 12694 33214 12794 33836
rect 12694 32886 12710 33214
rect 12782 32886 12794 33214
rect 12694 32870 12794 32886
rect 15821 27236 15920 38120
rect 12811 27137 15920 27236
rect 12811 26512 12910 27137
rect 12811 26080 12824 26512
rect 12898 26080 12910 26512
rect 12811 26067 12910 26080
rect 16120 20342 16220 43200
rect 16440 43140 16620 43160
rect 16440 43000 16460 43140
rect 16600 43000 16620 43140
rect 16440 42980 16620 43000
rect 12694 20242 16220 20342
rect 16480 20382 16580 42980
rect 16860 27300 16960 43400
rect 17140 34040 17240 43800
rect 17440 39824 17540 44260
rect 17440 39724 25516 39824
rect 25416 39258 25516 39724
rect 25416 38862 25432 39258
rect 25502 38862 25516 39258
rect 25416 38844 25516 38862
rect 17140 33940 25422 34040
rect 25322 33132 25422 33940
rect 25322 32804 25336 33132
rect 25408 32804 25422 33132
rect 25322 32792 25422 32804
rect 16860 27200 25602 27300
rect 16860 27174 16960 27200
rect 25502 26382 25602 27200
rect 25502 25988 25518 26382
rect 25586 25988 25602 26382
rect 25502 25970 25602 25988
rect 16480 20282 25938 20382
rect 12694 19464 12794 20242
rect 12694 19126 12706 19464
rect 12780 19126 12794 19464
rect 12694 19108 12794 19126
rect 25838 19334 25938 20282
rect 25838 18942 25852 19334
rect 25926 18942 25938 19334
rect 25838 18928 25938 18942
<< via2 >>
rect 14980 44480 15120 44600
rect 17400 44280 17580 44400
rect 15400 44040 15580 44200
rect 12656 38710 12734 39108
rect 17100 43820 17300 44000
rect 15780 43620 15960 43780
rect 16840 43420 16980 43540
rect 16100 43220 16240 43340
rect 12710 32886 12782 33214
rect 12824 26080 12898 26512
rect 16460 43000 16600 43140
rect 25432 38862 25502 39258
rect 25336 32804 25408 33132
rect 25518 25988 25586 26382
rect 12706 19126 12780 19464
rect 25852 18942 25926 19334
<< metal3 >>
rect 14960 44600 15140 44620
rect 14960 44480 14980 44600
rect 15120 44588 15140 44600
rect 29460 44600 29600 44620
rect 29460 44588 29480 44600
rect 15120 44495 29480 44588
rect 15120 44480 15140 44495
rect 14960 44460 15140 44480
rect 29460 44480 29480 44495
rect 29580 44480 29600 44600
rect 29460 44460 29600 44480
rect 17380 44400 17600 44420
rect 17380 44280 17400 44400
rect 17580 44386 17600 44400
rect 28720 44400 28880 44420
rect 28720 44386 28740 44400
rect 17580 44292 28740 44386
rect 17580 44280 17600 44292
rect 17380 44260 17600 44280
rect 28720 44280 28740 44292
rect 28860 44280 28880 44400
rect 28720 44260 28880 44280
rect 15380 44200 15600 44220
rect 15380 44040 15400 44200
rect 15580 44182 15600 44200
rect 27980 44200 28140 44220
rect 27980 44182 28000 44200
rect 15580 44088 28000 44182
rect 15580 44040 15600 44088
rect 15380 44020 15600 44040
rect 27980 44040 28000 44088
rect 28120 44040 28140 44200
rect 27980 44020 28140 44040
rect 17080 44000 17320 44020
rect 17080 43820 17100 44000
rect 17300 43956 17320 44000
rect 27220 44000 27420 44020
rect 27220 43956 27240 44000
rect 17300 43862 27240 43956
rect 17300 43820 17320 43862
rect 17080 43800 17320 43820
rect 27220 43820 27240 43862
rect 27400 43820 27420 44000
rect 27220 43800 27420 43820
rect 15760 43780 15980 43800
rect 15760 43620 15780 43780
rect 15960 43728 15980 43780
rect 26500 43760 26680 43780
rect 26500 43728 26520 43760
rect 15960 43634 26520 43728
rect 15960 43620 15980 43634
rect 15760 43600 15980 43620
rect 26500 43620 26520 43634
rect 26660 43620 26680 43760
rect 26500 43600 26680 43620
rect 16820 43540 17000 43560
rect 16820 43420 16840 43540
rect 16980 43524 17000 43540
rect 25720 43540 25960 43560
rect 25720 43524 25760 43540
rect 16980 43430 25760 43524
rect 16980 43420 17000 43430
rect 16820 43400 17000 43420
rect 25720 43420 25760 43430
rect 25940 43420 25960 43540
rect 25720 43400 25960 43420
rect 16080 43340 16260 43360
rect 16080 43220 16100 43340
rect 16240 43320 16260 43340
rect 25000 43340 25220 43360
rect 25000 43320 25020 43340
rect 16240 43226 25020 43320
rect 16240 43220 16260 43226
rect 16080 43200 16260 43220
rect 25000 43220 25020 43226
rect 25200 43220 25220 43340
rect 25000 43200 25220 43220
rect 16440 43140 16620 43160
rect 16440 43000 16460 43140
rect 16600 43128 16620 43140
rect 24260 43140 24480 43160
rect 24260 43128 24280 43140
rect 16600 43034 24280 43128
rect 16600 43000 16620 43034
rect 16440 42980 16620 43000
rect 24260 43000 24280 43034
rect 24460 43000 24480 43140
rect 24260 42980 24480 43000
rect 29335 39269 29658 39272
rect 2490 38596 5462 39012
rect 13930 38800 18246 39120
rect 26745 38951 29658 39269
rect 2490 2600 2906 38596
rect 29335 34518 29658 38951
rect 5090 34198 29658 34518
rect 5092 32668 5519 34198
rect 29335 34197 29658 34198
rect 5094 32368 5406 32668
rect 14054 32654 18248 32994
rect 26708 32836 29522 33156
rect 29204 28398 29520 32836
rect 5290 28082 29520 28398
rect 5296 25874 5636 28082
rect 14096 25960 18366 26280
rect 26804 25946 29360 26266
rect 5172 21674 5512 21690
rect 29040 21674 29360 25946
rect 5172 21354 29360 21674
rect 5172 18864 5512 21354
rect 13972 19136 18688 19456
rect 27154 19032 29640 19352
rect 2490 2500 2506 2600
rect 2888 2500 2906 2600
rect 2490 2396 2906 2500
rect 29325 1442 29636 19032
rect 26876 1430 29636 1442
rect 26876 1146 26910 1430
rect 27002 1146 29636 1430
rect 26876 1131 29636 1146
<< via3 >>
rect 29480 44480 29580 44600
rect 28740 44280 28860 44400
rect 28000 44040 28120 44200
rect 27240 43820 27400 44000
rect 26520 43620 26660 43760
rect 25760 43420 25940 43540
rect 25020 43220 25200 43340
rect 24280 43000 24460 43140
rect 2506 2500 2888 2600
rect 26910 1146 27002 1430
<< metal4 >>
rect 798 44486 858 45152
rect 1534 44486 1594 45152
rect 2270 44486 2330 45152
rect 3006 44486 3066 45152
rect 3742 44486 3802 45152
rect 4478 44486 4538 45152
rect 5214 44486 5274 45152
rect 5950 44486 6010 45152
rect 6686 44486 6746 45152
rect 7422 44486 7482 45152
rect 8158 44486 8218 45152
rect 8894 44486 8954 45152
rect 9630 44486 9690 45152
rect 10366 44486 10426 45152
rect 11102 44486 11162 45152
rect 11838 44486 11898 45152
rect 12574 44486 12634 45152
rect 13310 44486 13370 45152
rect 14046 44486 14106 45152
rect 14782 44486 14842 45152
rect 15518 44486 15578 45152
rect 16254 44486 16314 45152
rect 16990 44486 17050 45152
rect 17726 44486 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 798 44426 23156 44486
rect 1000 38600 1300 44152
rect 23096 42192 23156 44426
rect 24350 43160 24410 45152
rect 25086 43360 25146 45152
rect 25822 43560 25882 45152
rect 26558 43780 26618 45152
rect 27294 44020 27354 45152
rect 28030 44220 28090 45152
rect 28766 44420 28826 45152
rect 29502 44620 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 29460 44600 29600 44620
rect 29460 44480 29480 44600
rect 29580 44480 29600 44600
rect 29460 44460 29600 44480
rect 28720 44400 28880 44420
rect 28720 44280 28740 44400
rect 28860 44280 28880 44400
rect 28720 44260 28880 44280
rect 27980 44200 28140 44220
rect 27980 44040 28000 44200
rect 28120 44040 28140 44200
rect 27980 44020 28140 44040
rect 27220 44000 27420 44020
rect 27220 43820 27240 44000
rect 27400 43820 27420 44000
rect 27220 43800 27420 43820
rect 26500 43760 26680 43780
rect 26500 43620 26520 43760
rect 26660 43620 26680 43760
rect 26500 43600 26680 43620
rect 25720 43540 25960 43560
rect 25720 43420 25760 43540
rect 25940 43420 25960 43540
rect 25720 43400 25960 43420
rect 25000 43340 25220 43360
rect 25000 43220 25020 43340
rect 25200 43220 25220 43340
rect 25000 43200 25220 43220
rect 24260 43140 24480 43160
rect 24260 43000 24280 43140
rect 24460 43000 24480 43140
rect 24260 42980 24480 43000
rect 31506 42192 31806 44152
rect 23096 42132 31806 42192
rect 1000 37000 28800 38600
rect 1000 32600 1300 37000
rect 31506 36400 31806 42132
rect 5400 35000 31806 36400
rect 1000 31000 28800 32600
rect 1000 25600 1300 31000
rect 31506 30400 31806 35000
rect 5400 29000 31806 30400
rect 1000 24000 28800 25600
rect 1000 18400 1300 24000
rect 31506 23600 31806 29000
rect 5400 22200 31806 23600
rect 1000 17200 28800 18400
rect 1000 1000 1300 17200
rect 31506 16800 31806 22200
rect 5400 15400 31806 16800
rect 2417 2600 28525 2609
rect 2417 2500 2506 2600
rect 2888 2500 28525 2600
rect 2417 2491 28525 2500
rect 26896 1430 27016 1456
rect 26896 1146 26910 1430
rect 27002 1146 27016 1430
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 200
rect 13648 0 13768 200
rect 18064 0 18184 200
rect 22480 0 22600 200
rect 26896 0 27016 1146
rect 28407 482 28525 2491
rect 31506 1000 31806 15400
rect 28406 362 31432 482
rect 31312 0 31432 362
use bufferUnit  bufferUnit_0
timestamp 1713492510
transform 1 0 5996 0 1 34878
box -840 -120 9200 4280
use distortionUnit  distortionUnit_0
timestamp 1713492510
transform 1 0 6012 0 1 15202
box -840 -260 9200 4280
use distortionUnit  distortionUnit_2
timestamp 1713492510
transform 1 0 18784 0 1 34996
box -840 -260 9200 4280
use distortionUnit  distortionUnit_3
timestamp 1713492510
transform 1 0 6016 0 1 28952
box -840 -260 9200 4280
use distortionUnit  distortionUnit_4
timestamp 1713492510
transform 1 0 18748 0 1 28876
box -840 -260 9200 4280
use distortionUnit  distortionUnit_5
timestamp 1713492510
transform 1 0 6136 0 1 22248
box -840 -260 9200 4280
use distortionUnit  distortionUnit_6
timestamp 1713492510
transform 1 0 18844 0 1 22118
box -840 -260 9200 4280
use distortionUnit  distortionUnit_7
timestamp 1713492510
transform 1 0 19194 0 1 15072
box -840 -260 9200 4280
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 31506 1000 31806 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 1000 1000 1300 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
