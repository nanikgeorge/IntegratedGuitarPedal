magic
tech sky130A
magscale 1 2
timestamp 1713321159
<< nmos >>
rect -358 -73 -158 11
rect -100 -73 100 11
rect 158 -73 358 11
<< ndiff >>
rect -416 -1 -358 11
rect -416 -61 -404 -1
rect -370 -61 -358 -1
rect -416 -73 -358 -61
rect -158 -1 -100 11
rect -158 -61 -146 -1
rect -112 -61 -100 -1
rect -158 -73 -100 -61
rect 100 -1 158 11
rect 100 -61 112 -1
rect 146 -61 158 -1
rect 100 -73 158 -61
rect 358 -1 416 11
rect 358 -61 370 -1
rect 404 -61 416 -1
rect 358 -73 416 -61
<< ndiffc >>
rect -404 -61 -370 -1
rect -146 -61 -112 -1
rect 112 -61 146 -1
rect 370 -61 404 -1
<< poly >>
rect -358 83 -158 99
rect -358 49 -342 83
rect -174 49 -158 83
rect -358 11 -158 49
rect -100 83 100 99
rect -100 49 -84 83
rect 84 49 100 83
rect -100 11 100 49
rect 158 83 358 99
rect 158 49 174 83
rect 342 49 358 83
rect 158 11 358 49
rect -358 -99 -158 -73
rect -100 -99 100 -73
rect 158 -99 358 -73
<< polycont >>
rect -342 49 -174 83
rect -84 49 84 83
rect 174 49 342 83
<< locali >>
rect -358 49 -342 83
rect -174 49 -158 83
rect -100 49 -84 83
rect 84 49 100 83
rect 158 49 174 83
rect 342 49 358 83
rect -404 -1 -370 15
rect -404 -77 -370 -61
rect -146 -1 -112 15
rect -146 -77 -112 -61
rect 112 -1 146 15
rect 112 -77 146 -61
rect 370 -1 404 15
rect 370 -77 404 -61
<< viali >>
rect -342 49 -174 83
rect -84 49 84 83
rect 174 49 342 83
rect -404 -61 -370 -1
rect -146 -61 -112 -1
rect 112 -61 146 -1
rect 370 -61 404 -1
<< metal1 >>
rect -354 83 -162 89
rect -354 49 -342 83
rect -174 49 -162 83
rect -354 43 -162 49
rect -96 83 96 89
rect -96 49 -84 83
rect 84 49 96 83
rect -96 43 96 49
rect 162 83 354 89
rect 162 49 174 83
rect 342 49 354 83
rect 162 43 354 49
rect -410 -1 -364 11
rect -410 -61 -404 -1
rect -370 -61 -364 -1
rect -410 -73 -364 -61
rect -152 -1 -106 11
rect -152 -61 -146 -1
rect -112 -61 -106 -1
rect -152 -73 -106 -61
rect 106 -1 152 11
rect 106 -61 112 -1
rect 146 -61 152 -1
rect 106 -73 152 -61
rect 364 -1 410 11
rect 364 -61 370 -1
rect 404 -61 410 -1
rect 364 -73 410 -61
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.42 l 1 m 1 nf 3 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
