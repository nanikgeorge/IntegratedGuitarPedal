* NGSPICE file created from distortionUnit_lowR.ext - technology: sky130A

.subckt distortion_unit VDD CTRL IN OUT VSS
X0 a_1740_1605# a_1740_1605# VDD.t38 VDD.t37 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1 VDD.t36 a_1740_1605# tgate_1.IN VDD.t35 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2 tgate_1.IN a_1740_1605# VDD.t34 VDD.t33 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3 a_1740_1605# IN.t4 a_1998_1605# VSS.t29 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X4 a_1998_1605# IN.t5 a_1740_1605# VSS.t27 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X5 tgate_1.CTRLB CTRL.t0 VDD.t16 sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VSS.t38 a_896_1150# a_1998_1605# VSS.t37 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X7 VDD.t17 CTRL.t1 tgate_1.CTRLB sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8 a_1998_1605# a_896_1150# VSS.t36 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X9 VDD.t13 CTRL.t2 tgate_1.CTRLB sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VDD a_896_1150# VSS sky130_fd_pr__res_xhigh_po_0p35 l=26.11
X11 VSS.t34 a_896_1150# a_896_1150# VSS.t33 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X12 tgate_1.CTRLB CTRL.t3 VDD.t10 sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 tgate_1.CTRLB CTRL.t4 VDD.t6 sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X14 tgate_1.CTRLB CTRL.t5 VSS.t46 VSS.t45 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VDD.t32 a_1740_1605# a_1740_1605# VDD.t31 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X16 tgate_1.IN tgate_1.CTRLB OUT.t1 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X17 a_1740_1605# VDD.t3 VDD.t5 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X18 VDD.t30 a_1740_1605# a_1740_1605# VDD.t29 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X19 VDD.t11 CTRL.t6 tgate_1.CTRLB sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 a_1740_1605# IN.t6 a_1998_1605# VSS.t37 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X21 VSS.t24 VSS.t22 VSS.t24 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X22 OUT.t5 CTRL.t7 tgate_1.IN VSS.t53 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X23 VSS.t59 CTRL.t8 tgate_1.CTRLB VSS.t58 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 OUT.t7 CTRL.t9 IN.t3 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X25 a_1998_1605# myOpamp_0.INn tgate_1.IN VSS.t35 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X26 VSS.t21 VSS.t19 VSS.t20 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0 ps=0 w=0.42 l=1
X27 VSS.t18 VSS.t16 VSS.t18 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X28 tgate_1.IN myOpamp_0.INn a_1998_1605# VSS.t33 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X29 IN.t1 tgate_1.CTRLB OUT.t3 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X30 VDD.t12 a_896_1150# VSS.t49 sky130_fd_pr__res_xhigh_po_0p35 l=0.16
X31 VSS myOpamp_0.INn VSS.t39 sky130_fd_pr__res_xhigh_po_0p69 l=4
X32 tgate_1.CTRLB CTRL.t10 VSS.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X33 tgate_1.IN myOpamp_0.INn VSS.t44 sky130_fd_pr__res_xhigh_po_0p69 l=10
X34 VDD.t28 a_1740_1605# tgate_1.IN VDD.t27 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X35 VDD.t2 VDD.t0 tgate_1.IN VDD.t1 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X36 tgate_1.CTRLB CTRL.t11 VSS.t57 VSS.t56 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X37 tgate_1.IN a_1740_1605# VDD.t26 VDD.t25 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X38 tgate_1.IN a_1740_1605# VDD.t22 VDD.t21 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X39 a_1740_1605# VSS.t13 VSS.t15 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X40 a_1998_1605# IN.t7 a_1740_1605# VSS.t23 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X41 a_1998_1605# IN.t8 a_1740_1605# VSS.t17 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X42 a_1998_1605# a_896_1150# VSS.t32 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X43 VSS.t12 VSS.t11 VSS.t12 VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X44 tgate_1.CTRLB CTRL.t12 VDD.t15 sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X45 VSS.t10 VSS.t8 VSS.t10 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X46 VSS.t7 VSS.t5 VSS.t7 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X47 OUT.t0 tgate_1.CTRLB tgate_1.IN VDD.t7 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X48 tgate_1.CTRLB CTRL.t13 VSS.t55 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X49 a_1740_1605# a_1740_1605# VDD.t24 VDD.t23 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X50 VDD.t20 a_1740_1605# a_1740_1605# VDD.t19 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X51 tgate_1.IN CTRL.t14 OUT.t4 VSS.t50 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X52 VSS.t52 CTRL.t15 tgate_1.CTRLB VSS.t51 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X53 a_1998_1605# myOpamp_0.INn tgate_1.IN VSS.t31 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X54 VSS.t4 VSS.t2 tgate_1.IN VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X55 VSS.t30 a_896_1150# a_1998_1605# VSS.t29 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X56 a_896_1150# a_896_1150# VSS.t28 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X57 tgate_1.IN myOpamp_0.INn a_1998_1605# VSS.t9 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X58 tgate_1.IN myOpamp_0.INn a_1998_1605# VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X59 IN.t2 CTRL.t16 OUT.t6 VDD.t9 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X60 VDD.t18 CTRL.t17 tgate_1.CTRLB sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X61 VSS.t43 CTRL.t18 tgate_1.CTRLB VSS.t42 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X62 OUT.t2 tgate_1.CTRLB IN.t0 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X63 VSS.t48 CTRL.t19 tgate_1.CTRLB VSS.t47 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
R0 VDD.n14 VDD.n13 18810
R1 VDD.n15 VDD.n14 18786.2
R2 VDD.n15 VDD.n6 18786.2
R3 VDD.n13 VDD.n6 18667.5
R4 VDD.n16 VDD.n4 7334.54
R5 VDD.n12 VDD.n5 7332.73
R6 VDD.n16 VDD.n5 7312.73
R7 VDD.n12 VDD.n4 7300
R8 VDD.n41 VDD.n39 4136.47
R9 VDD.n48 VDD.n46 4136.47
R10 VDD.n41 VDD.n38 2068.24
R11 VDD.n48 VDD.n45 2068.24
R12 VDD.n10 VDD.n8 781.188
R13 VDD.n18 VDD.n2 779.442
R14 VDD.n17 VDD.n3 779.056
R15 VDD.n11 VDD.n7 778.668
R16 VDD.t21 VDD.t1 478.712
R17 VDD.t29 VDD.t21 478.712
R18 VDD.t37 VDD.t29 478.712
R19 VDD.t35 VDD.t37 478.712
R20 VDD.t33 VDD.t35 478.712
R21 VDD.t19 VDD.t23 478.712
R22 VDD.t23 VDD.t27 478.712
R23 VDD.t27 VDD.t25 478.712
R24 VDD.t25 VDD.t31 478.712
R25 VDD.t31 VDD.t4 478.712
R26 VDD.n41 VDD.t9 452.676
R27 VDD.t14 VDD.n39 452.676
R28 VDD.n48 VDD.t8 452.676
R29 VDD.t7 VDD.n46 452.676
R30 VDD.n67 VDD.t6 342.377
R31 VDD.n57 VDD.t17 338.892
R32 VDD.n72 VDD.n65 320.976
R33 VDD.n64 VDD.n54 320.976
R34 VDD.n62 VDD.n55 320.976
R35 VDD.n32 VDD.t12 269.151
R36 VDD.n31 VDD.t19 269.043
R37 VDD.n26 VDD.t5 228.215
R38 VDD.n21 VDD.t2 228.215
R39 VDD.t9 VDD.n40 215.757
R40 VDD.n40 VDD.t14 215.757
R41 VDD.t8 VDD.n47 215.757
R42 VDD.n47 VDD.t7 215.757
R43 VDD.n31 VDD.t33 209.668
R44 VDD.n28 VDD.n27 199.851
R45 VDD.n30 VDD.n29 199.851
R46 VDD.n23 VDD.n22 199.851
R47 VDD.n25 VDD.n24 199.851
R48 VDD.n35 VDD.n34 199.851
R49 VDD.n39 VDD.n37 163.684
R50 VDD.n46 VDD.n44 163.684
R51 VDD.n21 VDD.t0 120.855
R52 VDD.n26 VDD.t3 120.749
R53 VDD.n42 VDD.n37 113.915
R54 VDD.n49 VDD.n44 113.915
R55 VDD.n42 VDD.n41 47.0382
R56 VDD.n49 VDD.n48 47.0382
R57 VDD.n32 VDD.n31 38.8096
R58 VDD.n57 VDD 35.5709
R59 VDD.n61 VDD.n56 34.6358
R60 VDD.n74 VDD.n73 34.6358
R61 VDD.n71 VDD.n66 34.6358
R62 VDD.n64 VDD.n63 32.0005
R63 VDD.n63 VDD.n62 31.2476
R64 VDD.n27 VDD.t26 28.5655
R65 VDD.n27 VDD.t32 28.5655
R66 VDD.n29 VDD.t24 28.5655
R67 VDD.n29 VDD.t28 28.5655
R68 VDD.n22 VDD.t22 28.5655
R69 VDD.n22 VDD.t30 28.5655
R70 VDD.n24 VDD.t38 28.5655
R71 VDD.n24 VDD.t36 28.5655
R72 VDD.n34 VDD.t34 28.5655
R73 VDD.n34 VDD.t20 28.5655
R74 VDD.n65 VDD.t16 26.5955
R75 VDD.n65 VDD.t13 26.5955
R76 VDD.n54 VDD.t15 26.5955
R77 VDD.n54 VDD.t18 26.5955
R78 VDD.n55 VDD.t10 26.5955
R79 VDD.n55 VDD.t11 26.5955
R80 VDD.n73 VDD.n72 25.977
R81 VDD.n40 VDD.n38 20.5561
R82 VDD.n47 VDD.n45 20.5561
R83 VDD.n57 VDD.n56 18.824
R84 VDD.n38 VDD.n37 18.7435
R85 VDD.n45 VDD.n44 18.7435
R86 VDD.n67 VDD.n66 13.5534
R87 VDD VDD.n42 11.4981
R88 VDD VDD.n49 11.4981
R89 VDD.n68 VDD.n67 11.1829
R90 VDD.n58 VDD.n57 9.3005
R91 VDD.n59 VDD.n56 9.3005
R92 VDD.n61 VDD.n60 9.3005
R93 VDD.n63 VDD.n52 9.3005
R94 VDD.n75 VDD.n74 9.3005
R95 VDD.n73 VDD.n53 9.3005
R96 VDD.n71 VDD.n70 9.3005
R97 VDD.n69 VDD.n66 9.3005
R98 VDD.n72 VDD.n71 8.65932
R99 VDD.n8 VDD.n5 5.0005
R100 VDD.n14 VDD.n5 5.0005
R101 VDD.n7 VDD.n4 4.86892
R102 VDD.n6 VDD.n4 4.86892
R103 VDD.n62 VDD.n61 3.38874
R104 VDD.n51 VDD.n50 3.28283
R105 VDD.n51 VDD.n43 3.19667
R106 VDD.n74 VDD.n64 2.63579
R107 VDD.n19 VDD.n1 2.4755
R108 VDD.n9 VDD.n1 2.4755
R109 VDD.n9 VDD.n0 2.463
R110 VDD.n17 VDD.n16 2.34227
R111 VDD.n16 VDD.n15 2.34227
R112 VDD.n12 VDD.n11 2.34227
R113 VDD.n13 VDD.n12 2.34227
R114 VDD.n20 VDD.n0 2.10363
R115 VDD.n18 VDD.n17 1.93989
R116 VDD.n77 VDD.n76 1.02714
R117 VDD.n7 VDD.n2 0.970197
R118 VDD.n11 VDD.n10 0.970197
R119 VDD.n8 VDD.n3 0.970197
R120 VDD.n23 VDD.n21 0.890989
R121 VDD.n28 VDD.n26 0.760446
R122 VDD.n77 VDD.n51 0.419651
R123 VDD.n30 VDD.n28 0.40675
R124 VDD.n25 VDD.n23 0.40675
R125 VDD.n35 VDD.n25 0.40675
R126 VDD.n20 VDD.n19 0.359875
R127 VDD.n3 VDD.n1 0.258833
R128 VDD.n2 VDD.n0 0.258833
R129 VDD.n78 VDD.n77 0.257907
R130 VDD.n35 VDD.n33 0.208833
R131 VDD.n33 VDD.n30 0.188
R132 VDD.n33 VDD.n32 0.1865
R133 VDD.n78 VDD 0.15243
R134 VDD.n10 VDD.n9 0.121279
R135 VDD.n19 VDD.n18 0.121279
R136 VDD.n59 VDD.n58 0.120292
R137 VDD.n60 VDD.n59 0.120292
R138 VDD.n60 VDD.n52 0.120292
R139 VDD.n75 VDD.n53 0.120292
R140 VDD.n70 VDD.n53 0.120292
R141 VDD.n70 VDD.n69 0.120292
R142 VDD.n69 VDD.n68 0.120292
R143 VDD.n76 VDD.n75 0.115083
R144 VDD VDD.n80 0.096686
R145 VDD.n36 VDD.n35 0.0948367
R146 VDD.n36 VDD.n20 0.0691538
R147 VDD.n79 VDD.n36 0.0614341
R148 VDD.n58 VDD 0.0603958
R149 VDD VDD.n79 0.0562442
R150 VDD.n43 VDD 0.0459545
R151 VDD.n50 VDD 0.0459545
R152 VDD.n43 VDD 0.0338333
R153 VDD.n50 VDD 0.0338333
R154 VDD.n68 VDD 0.0226354
R155 VDD.n79 VDD.n78 0.00599114
R156 VDD.n76 VDD.n52 0.00570833
R157 IN.n4 IN.t2 223.565
R158 IN.n7 IN.t3 223.565
R159 IN.n0 IN.t8 118.769
R160 IN.n3 IN.t7 118.621
R161 IN.n2 IN.t4 118.005
R162 IN.n1 IN.t5 118.005
R163 IN.n0 IN.t6 118.005
R164 IN.n6 IN.n5 90.2112
R165 IN.n6 IN.n4 66.2405
R166 IN.n7 IN.n6 63.2157
R167 IN.n5 IN.t0 17.4005
R168 IN.n5 IN.t1 17.4005
R169 IN.n8 IN.n4 5.54823
R170 IN.n8 IN.n7 5.18686
R171 IN.n9 IN 4.4438
R172 IN IN.n3 2.77717
R173 IN.n1 IN.n0 2.66195
R174 IN.n3 IN.n2 1.71868
R175 IN.n2 IN.n1 0.764886
R176 IN IN.n9 0.490406
R177 IN IN.n8 0.244818
R178 IN.n9 IN 0.0129412
R179 VSS.n29 VSS.n28 80785
R180 VSS.n66 VSS.n65 27500
R181 VSS.n66 VSS.t49 10325.8
R182 VSS.n78 VSS.n60 10285.8
R183 VSS.n67 VSS.n60 10253
R184 VSS.n78 VSS.n61 10250
R185 VSS.n67 VSS.n61 10187.3
R186 VSS.n27 VSS.n26 9815.24
R187 VSS.n30 VSS.n27 9815.24
R188 VSS.n26 VSS.n17 9815.24
R189 VSS.n30 VSS.n17 9815.24
R190 VSS.n96 VSS.n6 9562.45
R191 VSS.n28 VSS.t39 7047.59
R192 VSS.n100 VSS.n3 6732.76
R193 VSS.n94 VSS.t39 6660.69
R194 VSS.n90 VSS.n18 6338.76
R195 VSS.n22 VSS.n18 6338.76
R196 VSS.n90 VSS.n19 6338.76
R197 VSS.n22 VSS.n19 6338.76
R198 VSS.n92 VSS.n5 6309.89
R199 VSS.n6 VSS.n5 4126.19
R200 VSS.n100 VSS.n4 3366.38
R201 VSS.n95 VSS.n94 2126.67
R202 VSS.n9 VSS.n7 1683.19
R203 VSS.n14 VSS.n7 1683.19
R204 VSS.t51 VSS.n92 1511.05
R205 VSS.n65 VSS.t3 1302.55
R206 VSS.t25 VSS.n10 1198.65
R207 VSS.n15 VSS.t26 1198.65
R208 VSS.n99 VSS.t53 1053.4
R209 VSS.t50 VSS.n97 1053.4
R210 VSS.n96 VSS.n95 967.52
R211 VSS.n91 VSS.n17 862.333
R212 VSS.n12 VSS.n7 841.596
R213 VSS.t3 VSS.t6 803.966
R214 VSS.t6 VSS.t17 803.966
R215 VSS.t17 VSS.t37 803.966
R216 VSS.t37 VSS.t35 803.966
R217 VSS.t35 VSS.t33 803.966
R218 VSS.t27 VSS.t29 803.966
R219 VSS.t9 VSS.t31 803.966
R220 VSS.t23 VSS.t9 803.966
R221 VSS.t14 VSS.t23 803.966
R222 VSS VSS.t54 785.428
R223 VSS.t56 VSS.t51 673.225
R224 VSS.t58 VSS.t56 673.225
R225 VSS.t0 VSS.t58 673.225
R226 VSS.t47 VSS.t0 673.225
R227 VSS.t45 VSS.t47 673.225
R228 VSS.t42 VSS.t45 673.225
R229 VSS.t54 VSS.t42 673.225
R230 VSS.n71 VSS.n62 666.376
R231 VSS.n77 VSS.n76 665.019
R232 VSS.n70 VSS.n69 664.242
R233 VSS.n68 VSS.n63 661.915
R234 VSS.t49 VSS.t14 660.674
R235 VSS.n25 VSS.n24 637.741
R236 VSS.n25 VSS.n23 637.741
R237 VSS.n31 VSS.n23 637.741
R238 VSS.n11 VSS.t25 636.323
R239 VSS.n11 VSS.t26 636.323
R240 VSS.t29 VSS.n79 629.462
R241 VSS.t53 VSS.n98 559.212
R242 VSS.n98 VSS.t50 559.212
R243 VSS.n93 VSS 536.976
R244 VSS.n92 VSS 469.406
R245 VSS.n80 VSS.t33 414.449
R246 VSS.n87 VSS.n86 411.495
R247 VSS.n88 VSS.n87 398.683
R248 VSS.n80 VSS.t27 389.519
R249 VSS.n89 VSS.n20 347.647
R250 VSS.n32 VSS.n21 287.356
R251 VSS.n118 VSS.t55 287.151
R252 VSS.n107 VSS.t52 284.024
R253 VSS.n10 VSS.n6 261.435
R254 VSS.n96 VSS.n15 261.435
R255 VSS.n14 VSS.n13 254.685
R256 VSS.n52 VSS.t21 236.113
R257 VSS.t12 VSS.n36 235.764
R258 VSS.n3 VSS.n2 232.597
R259 VSS.n99 VSS.n5 229.755
R260 VSS.n97 VSS.n96 229.755
R261 VSS.n29 VSS.t44 218.202
R262 VSS.n112 VSS.n106 207.213
R263 VSS.n125 VSS.n113 207.213
R264 VSS.n115 VSS.n114 207.213
R265 VSS.n86 VSS.n22 199.829
R266 VSS.t44 VSS.n16 197.768
R267 VSS.n28 VSS.n22 195
R268 VSS.n27 VSS.n23 195
R269 VSS.t44 VSS.n27 195
R270 VSS.n90 VSS.n89 195
R271 VSS.n91 VSS.n90 195
R272 VSS.n24 VSS.n17 195
R273 VSS.n57 VSS.n56 194.805
R274 VSS.n43 VSS.n42 194.542
R275 VSS.n59 VSS.n58 194.463
R276 VSS.n45 VSS.n44 194.463
R277 VSS.n53 VSS.n52 194.3
R278 VSS.n55 VSS.n54 194.3
R279 VSS.n41 VSS.n40 194.3
R280 VSS.n38 VSS.n37 194.3
R281 VSS.n65 VSS.n60 189.166
R282 VSS.n79 VSS.t31 174.505
R283 VSS.n9 VSS.n8 147.038
R284 VSS.n101 VSS.n100 147.038
R285 VSS.n10 VSS.n9 146.25
R286 VSS.n15 VSS.n14 146.25
R287 VSS.n97 VSS.n3 146.25
R288 VSS.n100 VSS.n99 146.25
R289 VSS.n93 VSS.n91 143
R290 VSS.n49 VSS.t13 118.005
R291 VSS.n35 VSS.t2 118.005
R292 VSS.n86 VSS.n85 113.481
R293 VSS.n50 VSS.t19 104.028
R294 VSS.n48 VSS.t22 104.028
R295 VSS.n47 VSS.t8 104.028
R296 VSS.n33 VSS.t16 104.028
R297 VSS.n39 VSS.t5 104.028
R298 VSS.n34 VSS.t11 104.028
R299 VSS.n101 VSS.n2 92.9264
R300 VSS.n13 VSS.n8 88.4348
R301 VSS.n49 VSS.t15 87.6949
R302 VSS.n35 VSS.t4 87.5315
R303 VSS.n24 VSS.n21 80.224
R304 VSS.t49 VSS.n61 77.0353
R305 VSS.n32 VSS.n31 67.8728
R306 VSS.n13 VSS.n12 65.0005
R307 VSS.n12 VSS.n11 65.0005
R308 VSS.n98 VSS.n4 65.0005
R309 VSS.n4 VSS.n2 59.3637
R310 VSS.n94 VSS.n93 58.6672
R311 VSS.n95 VSS.n16 46.7261
R312 VSS.n56 VSS.t32 41.4291
R313 VSS.n56 VSS.t10 41.4291
R314 VSS.t24 VSS.n53 41.4291
R315 VSS.n53 VSS.t20 41.4291
R316 VSS.t10 VSS.n55 41.4291
R317 VSS.n55 VSS.t24 41.4291
R318 VSS.n58 VSS.t28 41.4291
R319 VSS.n58 VSS.t30 41.4291
R320 VSS.n42 VSS.t18 41.4291
R321 VSS.n42 VSS.t38 41.4291
R322 VSS.n41 VSS.t7 41.4291
R323 VSS.t18 VSS.n41 41.4291
R324 VSS.n37 VSS.t12 41.4291
R325 VSS.n37 VSS.t7 41.4291
R326 VSS.n44 VSS.t36 41.4291
R327 VSS.n44 VSS.t34 41.4291
R328 VSS.n85 VSS.n20 36.4805
R329 VSS VSS.n107 35.197
R330 VSS.n111 VSS.n110 34.6358
R331 VSS.n124 VSS.n123 34.6358
R332 VSS.n120 VSS.n119 34.6358
R333 VSS.n126 VSS.n125 32.0005
R334 VSS.n126 VSS.n112 31.2476
R335 VSS.n81 VSS.n80 26.2219
R336 VSS.n123 VSS.n115 25.977
R337 VSS.n106 VSS.t57 24.9236
R338 VSS.n106 VSS.t59 24.9236
R339 VSS.n113 VSS.t1 24.9236
R340 VSS.n113 VSS.t48 24.9236
R341 VSS.n114 VSS.t46 24.9236
R342 VSS.n114 VSS.t43 24.9236
R343 VSS.n87 VSS.n19 23.4005
R344 VSS.n19 VSS.t39 23.4005
R345 VSS.n20 VSS.n18 23.4005
R346 VSS.n18 VSS.t39 23.4005
R347 VSS.n63 VSS.n61 20.8934
R348 VSS.n70 VSS.n60 20.8934
R349 VSS.n110 VSS.n107 18.824
R350 VSS.n26 VSS.n16 17.511
R351 VSS.n31 VSS.n30 13.6052
R352 VSS.n30 VSS.n29 13.6052
R353 VSS.n26 VSS.n25 13.6052
R354 VSS.n119 VSS.n118 13.5534
R355 VSS.n89 VSS.n88 13.177
R356 VSS.n8 VSS 11.4981
R357 VSS VSS.n101 11.4981
R358 VSS.n118 VSS.n117 11.1829
R359 VSS.n108 VSS.n107 9.3005
R360 VSS.n110 VSS.n109 9.3005
R361 VSS.n111 VSS.n104 9.3005
R362 VSS.n127 VSS.n126 9.3005
R363 VSS.n124 VSS.n105 9.3005
R364 VSS.n123 VSS.n122 9.3005
R365 VSS.n121 VSS.n120 9.3005
R366 VSS.n119 VSS.n116 9.3005
R367 VSS.n120 VSS.n115 8.65932
R368 VSS.n68 VSS.n67 8.23994
R369 VSS.n67 VSS.n66 8.23994
R370 VSS.n78 VSS.n77 8.23994
R371 VSS.n79 VSS.n78 8.23994
R372 VSS.n88 VSS.n21 4.3205
R373 VSS.n103 VSS.n1 3.45067
R374 VSS.n112 VSS.n111 3.38874
R375 VSS.n103 VSS.n102 2.87883
R376 VSS.n125 VSS.n124 2.63579
R377 VSS.n84 VSS.n32 2.45057
R378 VSS.n75 VSS.n64 2.09737
R379 VSS.n75 VSS.n74 2.09737
R380 VSS.n72 VSS.n64 2.09113
R381 VSS.n69 VSS.n68 1.93989
R382 VSS.n73 VSS.n72 1.72862
R383 VSS.n129 VSS.n128 1.24162
R384 VSS.n76 VSS.n63 0.970197
R385 VSS.n77 VSS.n62 0.970197
R386 VSS.n71 VSS.n70 0.970197
R387 VSS.n59 VSS.n57 0.927299
R388 VSS.n85 VSS.n84 0.846456
R389 VSS.n45 VSS.n43 0.690273
R390 VSS.n129 VSS.n103 0.6315
R391 VSS.n57 VSS.n46 0.60675
R392 VSS.n57 VSS.n51 0.516045
R393 VSS.n47 VSS.n46 0.454213
R394 VSS.n74 VSS.n73 0.363
R395 VSS.n54 VSS.n46 0.347226
R396 VSS.n72 VSS.n71 0.344944
R397 VSS.n76 VSS.n75 0.344944
R398 VSS.n48 VSS.n47 0.319807
R399 VSS.n51 VSS.n50 0.291342
R400 VSS.n54 VSS.n51 0.22669
R401 VSS.n82 VSS.n45 0.216409
R402 VSS.n130 VSS.n129 0.212
R403 VSS.n81 VSS.n59 0.210727
R404 VSS.n84 VSS.n83 0.158833
R405 VSS.n52 VSS.n51 0.158238
R406 VSS.n130 VSS 0.14
R407 VSS.n69 VSS.n64 0.135283
R408 VSS.n74 VSS.n62 0.135283
R409 VSS.n109 VSS.n108 0.120292
R410 VSS.n109 VSS.n104 0.120292
R411 VSS.n127 VSS.n105 0.120292
R412 VSS.n122 VSS.n105 0.120292
R413 VSS.n122 VSS.n121 0.120292
R414 VSS.n121 VSS.n116 0.120292
R415 VSS.n117 VSS.n116 0.120292
R416 VSS.n128 VSS.n104 0.112479
R417 VSS.n83 VSS.n82 0.09425
R418 VSS VSS.n132 0.0899516
R419 VSS.n50 VSS.n49 0.0714406
R420 VSS.n108 VSS 0.0603958
R421 VSS.n131 VSS.n0 0.0584812
R422 VSS VSS.n131 0.0520484
R423 VSS VSS.n1 0.0459545
R424 VSS.n102 VSS 0.0459545
R425 VSS.n73 VSS.n0 0.0455
R426 VSS.n38 VSS.n34 0.0429342
R427 VSS.n39 VSS.n38 0.0429342
R428 VSS.n40 VSS.n39 0.0429342
R429 VSS.n40 VSS.n33 0.0429342
R430 VSS.n36 VSS.n35 0.0389615
R431 VSS.n43 VSS.n33 0.0340526
R432 VSS.n1 VSS 0.0338333
R433 VSS.n102 VSS 0.0338333
R434 VSS.n51 VSS.n48 0.0289653
R435 VSS.n117 VSS 0.0226354
R436 VSS.n128 VSS.n127 0.0083125
R437 VSS.n36 VSS.n34 0.00773684
R438 VSS.n82 VSS.n81 0.00618182
R439 VSS.n131 VSS.n130 0.00544203
R440 VSS.n83 VSS.n0 0.00154167
R441 CTRL.n1 CTRL.t1 212.081
R442 CTRL.n25 CTRL.t3 212.081
R443 CTRL.n23 CTRL.t6 212.081
R444 CTRL.n2 CTRL.t12 212.081
R445 CTRL.n18 CTRL.t17 212.081
R446 CTRL.n3 CTRL.t0 212.081
R447 CTRL.n13 CTRL.t2 212.081
R448 CTRL.n11 CTRL.t4 212.081
R449 CTRL.n12 CTRL 163.264
R450 CTRL.n15 CTRL.n14 152
R451 CTRL.n17 CTRL.n16 152
R452 CTRL.n20 CTRL.n19 152
R453 CTRL.n22 CTRL.n21 152
R454 CTRL.n24 CTRL.n0 152
R455 CTRL CTRL.n26 152
R456 CTRL.n1 CTRL.t15 139.78
R457 CTRL.n25 CTRL.t11 139.78
R458 CTRL.n23 CTRL.t8 139.78
R459 CTRL.n2 CTRL.t10 139.78
R460 CTRL.n18 CTRL.t19 139.78
R461 CTRL.n3 CTRL.t5 139.78
R462 CTRL.n13 CTRL.t18 139.78
R463 CTRL.n11 CTRL.t13 139.78
R464 CTRL.n4 CTRL.t16 120.23
R465 CTRL.n4 CTRL.t9 120.228
R466 CTRL.n7 CTRL.t7 118.061
R467 CTRL.n7 CTRL.t14 118.058
R468 CTRL.n26 CTRL.n1 30.6732
R469 CTRL.n26 CTRL.n25 30.6732
R470 CTRL.n25 CTRL.n24 30.6732
R471 CTRL.n24 CTRL.n23 30.6732
R472 CTRL.n23 CTRL.n22 30.6732
R473 CTRL.n22 CTRL.n2 30.6732
R474 CTRL.n19 CTRL.n2 30.6732
R475 CTRL.n19 CTRL.n18 30.6732
R476 CTRL.n18 CTRL.n17 30.6732
R477 CTRL.n17 CTRL.n3 30.6732
R478 CTRL.n14 CTRL.n3 30.6732
R479 CTRL.n14 CTRL.n13 30.6732
R480 CTRL.n13 CTRL.n12 30.6732
R481 CTRL.n12 CTRL.n11 30.6732
R482 CTRL CTRL.n0 21.5045
R483 CTRL.n21 CTRL 19.4565
R484 CTRL CTRL.n20 17.4085
R485 CTRL CTRL.n15 13.3125
R486 CTRL.n16 CTRL.n10 13.0565
R487 CTRL.n15 CTRL 10.2405
R488 CTRL.n16 CTRL 8.1925
R489 CTRL.n20 CTRL 6.1445
R490 CTRL.n21 CTRL 4.0965
R491 CTRL.n10 CTRL.n9 3.2054
R492 CTRL.n10 CTRL 2.3045
R493 CTRL CTRL.n0 2.0485
R494 CTRL.n8 CTRL.n7 0.528909
R495 CTRL.n5 CTRL.n4 0.506182
R496 CTRL.n6 CTRL.n5 0.42675
R497 CTRL.n9 CTRL.n6 0.342556
R498 CTRL.n9 CTRL.n8 0.3415
R499 CTRL.n5 CTRL 0.170955
R500 CTRL.n8 CTRL 0.148227
R501 CTRL.n6 CTRL 0.01225
R502 OUT.n3 OUT.n1 199.941
R503 OUT.n10 OUT.n9 199.941
R504 OUT.n2 OUT.t3 83.7234
R505 OUT.n4 OUT.t2 83.7234
R506 OUT.n11 OUT.t4 83.7234
R507 OUT.n8 OUT.t5 83.7234
R508 OUT.n1 OUT.t6 28.5655
R509 OUT.n1 OUT.t7 28.5655
R510 OUT.n9 OUT.t1 28.5655
R511 OUT.n9 OUT.t0 28.5655
R512 OUT.n7 OUT.n6 1.15259
R513 OUT.n6 OUT.n5 0.938152
R514 OUT.n2 OUT.n0 0.5005
R515 OUT.n5 OUT.n4 0.5005
R516 OUT.n12 OUT.n11 0.5005
R517 OUT.n8 OUT.n7 0.5005
R518 OUT.n4 OUT.n3 0.478385
R519 OUT.n3 OUT.n2 0.478385
R520 OUT.n10 OUT.n8 0.478385
R521 OUT.n11 OUT.n10 0.478385
R522 OUT.n5 OUT.n0 0.364136
R523 OUT.n12 OUT.n7 0.364136
R524 OUT.n0 OUT 0.244818
R525 OUT OUT.n12 0.244818
R526 OUT.n6 OUT 0.0137188
C0 tgate_1.CTRLB CTRL 2.30483f
C1 VDD a_1740_1605# 4.48135f
C2 VDD CTRL 4.33897f
C3 OUT sky130_fd_sc_hd__tap_2_0.VPB 4.57e-19
C4 VDD a_896_1150# 0.128286f
C5 OUT IN 1.3678f
C6 OUT myOpamp_0.INn 0.005273f
C7 a_1740_1605# tgate_1.IN 2.35765f
C8 CTRL tgate_1.IN 0.795971f
C9 tgate_1.CTRLB sky130_fd_sc_hd__tap_2_0.VPB 0.175567f
C10 tgate_1.CTRLB OUT 1.62697f
C11 a_896_1150# tgate_1.IN 0.001336f
C12 IN a_1998_1605# 0.763261f
C13 myOpamp_0.INn a_1998_1605# 1.23683f
C14 VDD sky130_fd_sc_hd__tap_2_0.VPB 0.274328f
C15 myOpamp_0.INn IN 0.503808f
C16 VDD OUT 2.99895f
C17 tgate_1.CTRLB IN 0.258603f
C18 tgate_1.CTRLB myOpamp_0.INn 9.98e-19
C19 VDD a_1998_1605# 0.154599f
C20 VDD IN 6.86266f
C21 VDD myOpamp_0.INn 0.48498f
C22 tgate_1.CTRLB VDD 4.18127f
C23 OUT tgate_1.IN 1.38344f
C24 a_896_1150# a_1740_1605# 0.27522f
C25 a_1998_1605# tgate_1.IN 0.662032f
C26 IN tgate_1.IN 0.820736f
C27 myOpamp_0.INn tgate_1.IN 1.8069f
C28 tgate_1.CTRLB tgate_1.IN 1.18066f
C29 VDD tgate_1.IN 5.23663f
C30 CTRL sky130_fd_sc_hd__tap_2_0.VPB 0.278876f
C31 OUT CTRL 1.87653f
C32 a_1740_1605# a_1998_1605# 1.57848f
C33 IN a_1740_1605# 3.11184f
C34 myOpamp_0.INn a_1740_1605# 0.849481f
C35 CTRL IN 1.30918f
C36 myOpamp_0.INn CTRL 0.254411f
C37 a_896_1150# a_1998_1605# 1.5318f
C38 IN a_896_1150# 0.198383f
C39 myOpamp_0.INn a_896_1150# 1.1307f
C40 OUT VSS 5.986651f
C41 IN VSS 11.175117f
C42 CTRL VSS 7.482566f
C43 VDD VSS 55.798176f
C44 tgate_1.CTRLB VSS 4.58366f
C45 a_896_1150# VSS 5.5616f
C46 a_1998_1605# VSS 1.65017f
C47 myOpamp_0.INn VSS 7.25239f
C48 tgate_1.IN VSS 2.47159f
C49 a_1740_1605# VSS 2.78479f
C50 sky130_fd_sc_hd__tap_2_0.VPB VSS 1.14309f
C51 OUT.n0 VSS 0.15064f
C52 OUT.t6 VSS 0.003712f
C53 OUT.t7 VSS 0.003712f
C54 OUT.n1 VSS 0.007689f
C55 OUT.t3 VSS 0.013418f
C56 OUT.n2 VSS 0.107926f
C57 OUT.n3 VSS 0.101076f
C58 OUT.t2 VSS 0.013275f
C59 OUT.n4 VSS 0.105508f
C60 OUT.n5 VSS 0.264386f
C61 OUT.n6 VSS 0.694965f
C62 OUT.n7 VSS 0.338431f
C63 OUT.t5 VSS 0.013275f
C64 OUT.n8 VSS 0.105508f
C65 OUT.t1 VSS 0.003712f
C66 OUT.t0 VSS 0.003712f
C67 OUT.n9 VSS 0.007689f
C68 OUT.n10 VSS 0.101076f
C69 OUT.t4 VSS 0.013418f
C70 OUT.n11 VSS 0.107926f
C71 OUT.n12 VSS 0.15064f
C72 CTRL.n0 VSS 0.005024f
C73 CTRL.t1 VSS 0.009174f
C74 CTRL.t15 VSS 0.005406f
C75 CTRL.n1 VSS 0.012365f
C76 CTRL.t3 VSS 0.009174f
C77 CTRL.t11 VSS 0.005406f
C78 CTRL.t6 VSS 0.009174f
C79 CTRL.t8 VSS 0.005406f
C80 CTRL.t12 VSS 0.009174f
C81 CTRL.t10 VSS 0.005406f
C82 CTRL.n2 VSS 0.01323f
C83 CTRL.t17 VSS 0.009174f
C84 CTRL.t19 VSS 0.005406f
C85 CTRL.t0 VSS 0.009174f
C86 CTRL.t5 VSS 0.005406f
C87 CTRL.n3 VSS 0.01323f
C88 CTRL.t16 VSS 0.102501f
C89 CTRL.t9 VSS 0.1025f
C90 CTRL.n4 VSS 0.565618f
C91 CTRL.n5 VSS 0.383326f
C92 CTRL.n6 VSS 1.06549f
C93 CTRL.t7 VSS 0.099823f
C94 CTRL.t14 VSS 0.099822f
C95 CTRL.n7 VSS 0.57775f
C96 CTRL.n8 VSS 0.379137f
C97 CTRL.n9 VSS 2.01491f
C98 CTRL.n10 VSS 0.308073f
C99 CTRL.t2 VSS 0.009174f
C100 CTRL.t18 VSS 0.005406f
C101 CTRL.t4 VSS 0.009174f
C102 CTRL.t13 VSS 0.005406f
C103 CTRL.n11 VSS 0.012365f
C104 CTRL.n12 VSS 0.006469f
C105 CTRL.n13 VSS 0.01323f
C106 CTRL.n14 VSS 0.006055f
C107 CTRL.n15 VSS 0.005024f
C108 CTRL.n16 VSS 0.004532f
C109 CTRL.n17 VSS 0.006055f
C110 CTRL.n18 VSS 0.01323f
C111 CTRL.n19 VSS 0.006055f
C112 CTRL.n20 VSS 0.005024f
C113 CTRL.n21 VSS 0.005024f
C114 CTRL.n22 VSS 0.006055f
C115 CTRL.n23 VSS 0.01323f
C116 CTRL.n24 VSS 0.006055f
C117 CTRL.n25 VSS 0.01323f
C118 CTRL.n26 VSS 0.006055f
C119 IN.t8 VSS 0.107729f
C120 IN.t6 VSS 0.107375f
C121 IN.n0 VSS 0.133f
C122 IN.t5 VSS 0.107375f
C123 IN.n1 VSS 0.078467f
C124 IN.t4 VSS 0.107375f
C125 IN.n2 VSS 0.068105f
C126 IN.t7 VSS 0.10765f
C127 IN.n3 VSS 0.18673f
C128 IN.t2 VSS 0.024658f
C129 IN.n4 VSS 0.095276f
C130 IN.t0 VSS 0.006818f
C131 IN.t1 VSS 0.006818f
C132 IN.n5 VSS 0.022125f
C133 IN.n6 VSS 0.134918f
C134 IN.t3 VSS 0.024658f
C135 IN.n7 VSS 0.071178f
C136 IN.n8 VSS 0.815587f
C137 IN.n9 VSS 3.13504f
C138 VDD.n0 VSS 0.684451f
C139 VDD.n1 VSS 0.741033f
C140 VDD.n2 VSS 0.121361f
C141 VDD.n3 VSS 0.121301f
C142 VDD.n4 VSS 0.242751f
C143 VDD.n5 VSS 0.242931f
C144 VDD.n6 VSS 0.737821f
C145 VDD.n7 VSS 0.121241f
C146 VDD.n8 VSS 0.121631f
C147 VDD.n9 VSS 0.725011f
C148 VDD.n10 VSS 0.120918f
C149 VDD.n11 VSS 0.120532f
C150 VDD.n12 VSS 0.241301f
C151 VDD.n13 VSS 0.724075f
C152 VDD.n14 VSS 0.740574f
C153 VDD.n15 VSS 0.725946f
C154 VDD.n16 VSS 0.241542f
C155 VDD.n17 VSS 0.12074f
C156 VDD.n18 VSS 0.1208f
C157 VDD.n19 VSS 0.415366f
C158 VDD.n20 VSS 0.774972f
C159 VDD.t0 VSS 0.042525f
C160 VDD.t2 VSS 0.00963f
C161 VDD.n21 VSS 0.055724f
C162 VDD.t22 VSS 0.002621f
C163 VDD.t30 VSS 0.002621f
C164 VDD.n22 VSS 0.00542f
C165 VDD.n23 VSS 0.107629f
C166 VDD.t38 VSS 0.002621f
C167 VDD.t36 VSS 0.002621f
C168 VDD.n24 VSS 0.00542f
C169 VDD.n25 VSS 0.09048f
C170 VDD.t3 VSS 0.042497f
C171 VDD.t5 VSS 0.00963f
C172 VDD.n26 VSS 0.09949f
C173 VDD.t26 VSS 0.002621f
C174 VDD.t32 VSS 0.002621f
C175 VDD.n27 VSS 0.00542f
C176 VDD.n28 VSS 0.131214f
C177 VDD.t24 VSS 0.002621f
C178 VDD.t28 VSS 0.002621f
C179 VDD.n29 VSS 0.00542f
C180 VDD.n30 VSS 0.079092f
C181 VDD.t1 VSS 0.149472f
C182 VDD.t21 VSS 0.119393f
C183 VDD.t29 VSS 0.119393f
C184 VDD.t37 VSS 0.119393f
C185 VDD.t35 VSS 0.119393f
C186 VDD.t33 VSS 0.085842f
C187 VDD.t4 VSS 0.149472f
C188 VDD.t31 VSS 0.119393f
C189 VDD.t25 VSS 0.119393f
C190 VDD.t27 VSS 0.119393f
C191 VDD.t23 VSS 0.119393f
C192 VDD.t19 VSS 0.093246f
C193 VDD.n31 VSS -0.070015f
C194 VDD.t12 VSS 0.100561f
C195 VDD.n32 VSS 0.154476f
C196 VDD.n33 VSS 0.020607f
C197 VDD.t34 VSS 0.002621f
C198 VDD.t20 VSS 0.002621f
C199 VDD.n34 VSS 0.00542f
C200 VDD.n35 VSS 0.088934f
C201 VDD.n36 VSS 3.16797f
C202 VDD.n37 VSS 0.031907f
C203 VDD.n38 VSS 0.018389f
C204 VDD.n39 VSS 0.131251f
C205 VDD.t14 VSS 0.104641f
C206 VDD.n40 VSS 0.066226f
C207 VDD.t9 VSS 0.104641f
C208 VDD.n41 VSS 0.108423f
C209 VDD.n42 VSS 0.056743f
C210 VDD.n43 VSS 0.250005f
C211 VDD.n44 VSS 0.031907f
C212 VDD.n45 VSS 0.018389f
C213 VDD.n46 VSS 0.131251f
C214 VDD.t7 VSS 0.104641f
C215 VDD.n47 VSS 0.066226f
C216 VDD.t8 VSS 0.104641f
C217 VDD.n48 VSS 0.108423f
C218 VDD.n49 VSS 0.056743f
C219 VDD.n50 VSS 0.253103f
C220 VDD.n51 VSS 0.423553f
C221 VDD.n52 VSS 0.004165f
C222 VDD.n53 VSS 0.007983f
C223 VDD.t15 VSS 0.00244f
C224 VDD.t18 VSS 0.00244f
C225 VDD.n54 VSS 0.005239f
C226 VDD.t10 VSS 0.00244f
C227 VDD.t11 VSS 0.00244f
C228 VDD.n55 VSS 0.005239f
C229 VDD.n56 VSS 0.002182f
C230 VDD.t17 VSS 0.009291f
C231 VDD.n57 VSS 0.013237f
C232 VDD.n58 VSS 0.005987f
C233 VDD.n59 VSS 0.007983f
C234 VDD.n60 VSS 0.007983f
C235 VDD.n61 VSS 0.001552f
C236 VDD.n62 VSS 0.005973f
C237 VDD.n63 VSS 0.002581f
C238 VDD.n64 VSS 0.005973f
C239 VDD.t16 VSS 0.00244f
C240 VDD.t13 VSS 0.00244f
C241 VDD.n65 VSS 0.005239f
C242 VDD.n66 VSS 0.001967f
C243 VDD.t6 VSS 0.009292f
C244 VDD.n67 VSS 0.01092f
C245 VDD.n68 VSS 0.00498f
C246 VDD.n69 VSS 0.007983f
C247 VDD.n70 VSS 0.007983f
C248 VDD.n71 VSS 0.001767f
C249 VDD.n72 VSS 0.005973f
C250 VDD.n73 VSS 0.002474f
C251 VDD.n74 VSS 0.001521f
C252 VDD.n75 VSS 0.007809f
C253 VDD.n76 VSS 0.320831f
C254 VDD.n77 VSS 4.09046f
C255 VDD.n78 VSS 2.91097f
C256 VDD.n79 VSS 1.55655f
C257 VDD.n80 VSS 0.730658f
.ends

