magic
tech sky130A
magscale 1 2
timestamp 1713223699
<< nmos >>
rect -100 -19 100 81
<< ndiff >>
rect -158 69 -100 81
rect -158 -7 -146 69
rect -112 -7 -100 69
rect -158 -19 -100 -7
rect 100 69 158 81
rect 100 -7 112 69
rect 146 -7 158 69
rect 100 -19 158 -7
<< ndiffc >>
rect -146 -7 -112 69
rect 112 -7 146 69
<< poly >>
rect -100 81 100 107
rect -100 -57 100 -19
rect -100 -91 -84 -57
rect 84 -91 100 -57
rect -100 -107 100 -91
<< polycont >>
rect -84 -91 84 -57
<< locali >>
rect -146 69 -112 85
rect -146 -23 -112 -7
rect 112 69 146 85
rect 112 -23 146 -7
rect -100 -91 -84 -57
rect 84 -91 100 -57
<< viali >>
rect -146 -7 -112 69
rect 112 -7 146 69
rect -84 -91 84 -57
<< metal1 >>
rect -152 69 -106 81
rect -152 -7 -146 69
rect -112 -7 -106 69
rect -152 -19 -106 -7
rect 106 69 152 81
rect 106 -7 112 69
rect 146 -7 152 69
rect 106 -19 152 -7
rect -96 -57 96 -51
rect -96 -91 -84 -57
rect 84 -91 96 -57
rect -96 -97 96 -91
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.5 l 1 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
