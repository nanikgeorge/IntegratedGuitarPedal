magic
tech sky130A
magscale 1 2
timestamp 1713484462
<< nwell >>
rect -380 2920 5320 3120
rect -380 520 -180 2920
rect 1446 1932 4672 2444
rect 5120 520 5320 2920
rect 6727 3085 7577 3653
rect -380 320 5320 520
rect 6727 1625 7577 2193
rect 6520 289 7608 610
<< pwell >>
rect -80 2620 5020 2820
rect -80 820 1410 2620
rect 1440 1050 4670 1220
rect 4820 820 5020 2620
rect -80 620 5020 820
rect 3460 -260 5424 142
rect 5500 -260 5902 2904
rect 6727 2527 7577 3085
rect 6727 1067 7577 1625
rect 6592 49 7366 231
rect 7389 66 7567 223
rect 6592 45 6621 49
rect 6587 11 6621 45
<< nmos >>
rect 1540 1605 1740 1805
rect 1798 1605 1998 1805
rect 2056 1605 2256 1805
rect 2314 1605 2514 1805
rect 2572 1605 2772 1805
rect 2830 1605 3030 1805
rect 3088 1605 3288 1805
rect 3346 1605 3546 1805
rect 3604 1605 3804 1805
rect 3862 1605 4062 1805
rect 4120 1605 4320 1805
rect 4378 1605 4578 1805
rect 1540 1285 1740 1369
rect 1798 1285 1998 1369
rect 2056 1285 2256 1369
rect 2314 1285 2514 1369
rect 2572 1285 2772 1369
rect 2830 1285 3030 1369
rect 3088 1285 3288 1369
rect 3346 1285 3546 1369
rect 3604 1285 3804 1369
rect 3862 1285 4062 1369
rect 4120 1285 4320 1369
rect 4378 1285 4578 1369
rect 6923 2737 7123 2937
rect 7181 2737 7381 2937
rect 6923 1277 7123 1477
rect 7181 1277 7381 1477
<< scnmos >>
rect 6670 75 6700 205
rect 6754 75 6784 205
rect 6838 75 6868 205
rect 6922 75 6952 205
rect 7006 75 7036 205
rect 7090 75 7120 205
rect 7174 75 7204 205
rect 7258 75 7288 205
<< pmos >>
rect 6923 3233 7123 3433
rect 7181 3233 7381 3433
rect 1540 2032 1740 2232
rect 1798 2032 1998 2232
rect 2056 2032 2256 2232
rect 2314 2032 2514 2232
rect 2572 2032 2772 2232
rect 2830 2032 3030 2232
rect 3088 2032 3288 2232
rect 3346 2032 3546 2232
rect 3604 2032 3804 2232
rect 3862 2032 4062 2232
rect 4120 2032 4320 2232
rect 4378 2032 4578 2232
rect 6923 1773 7123 1973
rect 7181 1773 7381 1973
<< scpmoshvt >>
rect 6670 325 6700 525
rect 6754 325 6784 525
rect 6838 325 6868 525
rect 6922 325 6952 525
rect 7006 325 7036 525
rect 7090 325 7120 525
rect 7174 325 7204 525
rect 7258 325 7288 525
<< ndiff >>
rect 1482 1793 1540 1805
rect 1482 1617 1494 1793
rect 1528 1617 1540 1793
rect 1482 1605 1540 1617
rect 1740 1793 1798 1805
rect 1740 1617 1752 1793
rect 1786 1617 1798 1793
rect 1740 1605 1798 1617
rect 1998 1793 2056 1805
rect 1998 1617 2010 1793
rect 2044 1617 2056 1793
rect 1998 1605 2056 1617
rect 2256 1793 2314 1805
rect 2256 1617 2268 1793
rect 2302 1617 2314 1793
rect 2256 1605 2314 1617
rect 2514 1793 2572 1805
rect 2514 1617 2526 1793
rect 2560 1617 2572 1793
rect 2514 1605 2572 1617
rect 2772 1793 2830 1805
rect 2772 1617 2784 1793
rect 2818 1617 2830 1793
rect 2772 1605 2830 1617
rect 3030 1793 3088 1805
rect 3030 1617 3042 1793
rect 3076 1617 3088 1793
rect 3030 1605 3088 1617
rect 3288 1793 3346 1805
rect 3288 1617 3300 1793
rect 3334 1617 3346 1793
rect 3288 1605 3346 1617
rect 3546 1793 3604 1805
rect 3546 1617 3558 1793
rect 3592 1617 3604 1793
rect 3546 1605 3604 1617
rect 3804 1793 3862 1805
rect 3804 1617 3816 1793
rect 3850 1617 3862 1793
rect 3804 1605 3862 1617
rect 4062 1793 4120 1805
rect 4062 1617 4074 1793
rect 4108 1617 4120 1793
rect 4062 1605 4120 1617
rect 4320 1793 4378 1805
rect 4320 1617 4332 1793
rect 4366 1617 4378 1793
rect 4320 1605 4378 1617
rect 4578 1793 4636 1805
rect 4578 1617 4590 1793
rect 4624 1617 4636 1793
rect 4578 1605 4636 1617
rect 1482 1357 1540 1369
rect 1482 1297 1494 1357
rect 1528 1297 1540 1357
rect 1482 1285 1540 1297
rect 1740 1357 1798 1369
rect 1740 1297 1752 1357
rect 1786 1297 1798 1357
rect 1740 1285 1798 1297
rect 1998 1357 2056 1369
rect 1998 1297 2010 1357
rect 2044 1297 2056 1357
rect 1998 1285 2056 1297
rect 2256 1357 2314 1369
rect 2256 1297 2268 1357
rect 2302 1297 2314 1357
rect 2256 1285 2314 1297
rect 2514 1357 2572 1369
rect 2514 1297 2526 1357
rect 2560 1297 2572 1357
rect 2514 1285 2572 1297
rect 2772 1357 2830 1369
rect 2772 1297 2784 1357
rect 2818 1297 2830 1357
rect 2772 1285 2830 1297
rect 3030 1357 3088 1369
rect 3030 1297 3042 1357
rect 3076 1297 3088 1357
rect 3030 1285 3088 1297
rect 3288 1357 3346 1369
rect 3288 1297 3300 1357
rect 3334 1297 3346 1357
rect 3288 1285 3346 1297
rect 3546 1357 3604 1369
rect 3546 1297 3558 1357
rect 3592 1297 3604 1357
rect 3546 1285 3604 1297
rect 3804 1357 3862 1369
rect 3804 1297 3816 1357
rect 3850 1297 3862 1357
rect 3804 1285 3862 1297
rect 4062 1357 4120 1369
rect 4062 1297 4074 1357
rect 4108 1297 4120 1357
rect 4062 1285 4120 1297
rect 4320 1357 4378 1369
rect 4320 1297 4332 1357
rect 4366 1297 4378 1357
rect 4320 1285 4378 1297
rect 4578 1357 4636 1369
rect 4578 1297 4590 1357
rect 4624 1297 4636 1357
rect 4578 1285 4636 1297
rect 6865 2925 6923 2937
rect 6865 2749 6877 2925
rect 6911 2749 6923 2925
rect 6865 2737 6923 2749
rect 7123 2925 7181 2937
rect 7123 2749 7135 2925
rect 7169 2749 7181 2925
rect 7123 2737 7181 2749
rect 7381 2925 7439 2937
rect 7381 2749 7393 2925
rect 7427 2749 7439 2925
rect 7381 2737 7439 2749
rect 6865 1465 6923 1477
rect 6865 1289 6877 1465
rect 6911 1289 6923 1465
rect 6865 1277 6923 1289
rect 7123 1465 7181 1477
rect 7123 1289 7135 1465
rect 7169 1289 7181 1465
rect 7123 1277 7181 1289
rect 7381 1465 7439 1477
rect 7381 1289 7393 1465
rect 7427 1289 7439 1465
rect 7381 1277 7439 1289
rect 6618 121 6670 205
rect 6618 87 6626 121
rect 6660 87 6670 121
rect 6618 75 6670 87
rect 6700 189 6754 205
rect 6700 155 6710 189
rect 6744 155 6754 189
rect 6700 121 6754 155
rect 6700 87 6710 121
rect 6744 87 6754 121
rect 6700 75 6754 87
rect 6784 121 6838 205
rect 6784 87 6794 121
rect 6828 87 6838 121
rect 6784 75 6838 87
rect 6868 189 6922 205
rect 6868 155 6878 189
rect 6912 155 6922 189
rect 6868 121 6922 155
rect 6868 87 6878 121
rect 6912 87 6922 121
rect 6868 75 6922 87
rect 6952 121 7006 205
rect 6952 87 6962 121
rect 6996 87 7006 121
rect 6952 75 7006 87
rect 7036 189 7090 205
rect 7036 155 7046 189
rect 7080 155 7090 189
rect 7036 121 7090 155
rect 7036 87 7046 121
rect 7080 87 7090 121
rect 7036 75 7090 87
rect 7120 121 7174 205
rect 7120 87 7130 121
rect 7164 87 7174 121
rect 7120 75 7174 87
rect 7204 189 7258 205
rect 7204 155 7214 189
rect 7248 155 7258 189
rect 7204 121 7258 155
rect 7204 87 7214 121
rect 7248 87 7258 121
rect 7204 75 7258 87
rect 7288 121 7340 205
rect 7288 87 7298 121
rect 7332 87 7340 121
rect 7288 75 7340 87
<< pdiff >>
rect 6865 3421 6923 3433
rect 6865 3245 6877 3421
rect 6911 3245 6923 3421
rect 6865 3233 6923 3245
rect 7123 3421 7181 3433
rect 7123 3245 7135 3421
rect 7169 3245 7181 3421
rect 7123 3233 7181 3245
rect 7381 3421 7439 3433
rect 7381 3245 7393 3421
rect 7427 3245 7439 3421
rect 7381 3233 7439 3245
rect 1482 2220 1540 2232
rect 1482 2044 1494 2220
rect 1528 2044 1540 2220
rect 1482 2032 1540 2044
rect 1740 2220 1798 2232
rect 1740 2044 1752 2220
rect 1786 2044 1798 2220
rect 1740 2032 1798 2044
rect 1998 2220 2056 2232
rect 1998 2044 2010 2220
rect 2044 2044 2056 2220
rect 1998 2032 2056 2044
rect 2256 2220 2314 2232
rect 2256 2044 2268 2220
rect 2302 2044 2314 2220
rect 2256 2032 2314 2044
rect 2514 2220 2572 2232
rect 2514 2044 2526 2220
rect 2560 2044 2572 2220
rect 2514 2032 2572 2044
rect 2772 2220 2830 2232
rect 2772 2044 2784 2220
rect 2818 2044 2830 2220
rect 2772 2032 2830 2044
rect 3030 2220 3088 2232
rect 3030 2044 3042 2220
rect 3076 2044 3088 2220
rect 3030 2032 3088 2044
rect 3288 2220 3346 2232
rect 3288 2044 3300 2220
rect 3334 2044 3346 2220
rect 3288 2032 3346 2044
rect 3546 2220 3604 2232
rect 3546 2044 3558 2220
rect 3592 2044 3604 2220
rect 3546 2032 3604 2044
rect 3804 2220 3862 2232
rect 3804 2044 3816 2220
rect 3850 2044 3862 2220
rect 3804 2032 3862 2044
rect 4062 2220 4120 2232
rect 4062 2044 4074 2220
rect 4108 2044 4120 2220
rect 4062 2032 4120 2044
rect 4320 2220 4378 2232
rect 4320 2044 4332 2220
rect 4366 2044 4378 2220
rect 4320 2032 4378 2044
rect 4578 2220 4636 2232
rect 4578 2044 4590 2220
rect 4624 2044 4636 2220
rect 4578 2032 4636 2044
rect 6865 1961 6923 1973
rect 6865 1785 6877 1961
rect 6911 1785 6923 1961
rect 6865 1773 6923 1785
rect 7123 1961 7181 1973
rect 7123 1785 7135 1961
rect 7169 1785 7181 1961
rect 7123 1773 7181 1785
rect 7381 1961 7439 1973
rect 7381 1785 7393 1961
rect 7427 1785 7439 1961
rect 7381 1773 7439 1785
rect 6618 513 6670 525
rect 6618 479 6626 513
rect 6660 479 6670 513
rect 6618 445 6670 479
rect 6618 411 6626 445
rect 6660 411 6670 445
rect 6618 325 6670 411
rect 6700 513 6754 525
rect 6700 479 6710 513
rect 6744 479 6754 513
rect 6700 445 6754 479
rect 6700 411 6710 445
rect 6744 411 6754 445
rect 6700 377 6754 411
rect 6700 343 6710 377
rect 6744 343 6754 377
rect 6700 325 6754 343
rect 6784 513 6838 525
rect 6784 479 6794 513
rect 6828 479 6838 513
rect 6784 445 6838 479
rect 6784 411 6794 445
rect 6828 411 6838 445
rect 6784 325 6838 411
rect 6868 513 6922 525
rect 6868 479 6878 513
rect 6912 479 6922 513
rect 6868 445 6922 479
rect 6868 411 6878 445
rect 6912 411 6922 445
rect 6868 377 6922 411
rect 6868 343 6878 377
rect 6912 343 6922 377
rect 6868 325 6922 343
rect 6952 513 7006 525
rect 6952 479 6962 513
rect 6996 479 7006 513
rect 6952 445 7006 479
rect 6952 411 6962 445
rect 6996 411 7006 445
rect 6952 325 7006 411
rect 7036 513 7090 525
rect 7036 479 7046 513
rect 7080 479 7090 513
rect 7036 445 7090 479
rect 7036 411 7046 445
rect 7080 411 7090 445
rect 7036 377 7090 411
rect 7036 343 7046 377
rect 7080 343 7090 377
rect 7036 325 7090 343
rect 7120 513 7174 525
rect 7120 479 7130 513
rect 7164 479 7174 513
rect 7120 445 7174 479
rect 7120 411 7130 445
rect 7164 411 7174 445
rect 7120 325 7174 411
rect 7204 513 7258 525
rect 7204 479 7214 513
rect 7248 479 7258 513
rect 7204 445 7258 479
rect 7204 411 7214 445
rect 7248 411 7258 445
rect 7204 377 7258 411
rect 7204 343 7214 377
rect 7248 343 7258 377
rect 7204 325 7258 343
rect 7288 513 7340 525
rect 7288 479 7298 513
rect 7332 479 7340 513
rect 7288 445 7340 479
rect 7288 411 7298 445
rect 7332 411 7340 445
rect 7288 325 7340 411
<< ndiffc >>
rect 1494 1617 1528 1793
rect 1752 1617 1786 1793
rect 2010 1617 2044 1793
rect 2268 1617 2302 1793
rect 2526 1617 2560 1793
rect 2784 1617 2818 1793
rect 3042 1617 3076 1793
rect 3300 1617 3334 1793
rect 3558 1617 3592 1793
rect 3816 1617 3850 1793
rect 4074 1617 4108 1793
rect 4332 1617 4366 1793
rect 4590 1617 4624 1793
rect 1494 1297 1528 1357
rect 1752 1297 1786 1357
rect 2010 1297 2044 1357
rect 2268 1297 2302 1357
rect 2526 1297 2560 1357
rect 2784 1297 2818 1357
rect 3042 1297 3076 1357
rect 3300 1297 3334 1357
rect 3558 1297 3592 1357
rect 3816 1297 3850 1357
rect 4074 1297 4108 1357
rect 4332 1297 4366 1357
rect 4590 1297 4624 1357
rect 6877 2749 6911 2925
rect 7135 2749 7169 2925
rect 7393 2749 7427 2925
rect 6877 1289 6911 1465
rect 7135 1289 7169 1465
rect 7393 1289 7427 1465
rect 6626 87 6660 121
rect 6710 155 6744 189
rect 6710 87 6744 121
rect 6794 87 6828 121
rect 6878 155 6912 189
rect 6878 87 6912 121
rect 6962 87 6996 121
rect 7046 155 7080 189
rect 7046 87 7080 121
rect 7130 87 7164 121
rect 7214 155 7248 189
rect 7214 87 7248 121
rect 7298 87 7332 121
<< pdiffc >>
rect 6877 3245 6911 3421
rect 7135 3245 7169 3421
rect 7393 3245 7427 3421
rect 1494 2044 1528 2220
rect 1752 2044 1786 2220
rect 2010 2044 2044 2220
rect 2268 2044 2302 2220
rect 2526 2044 2560 2220
rect 2784 2044 2818 2220
rect 3042 2044 3076 2220
rect 3300 2044 3334 2220
rect 3558 2044 3592 2220
rect 3816 2044 3850 2220
rect 4074 2044 4108 2220
rect 4332 2044 4366 2220
rect 4590 2044 4624 2220
rect 6877 1785 6911 1961
rect 7135 1785 7169 1961
rect 7393 1785 7427 1961
rect 6626 479 6660 513
rect 6626 411 6660 445
rect 6710 479 6744 513
rect 6710 411 6744 445
rect 6710 343 6744 377
rect 6794 479 6828 513
rect 6794 411 6828 445
rect 6878 479 6912 513
rect 6878 411 6912 445
rect 6878 343 6912 377
rect 6962 479 6996 513
rect 6962 411 6996 445
rect 7046 479 7080 513
rect 7046 411 7080 445
rect 7046 343 7080 377
rect 7130 479 7164 513
rect 7130 411 7164 445
rect 7214 479 7248 513
rect 7214 411 7248 445
rect 7214 343 7248 377
rect 7298 479 7332 513
rect 7298 411 7332 445
<< psubdiff >>
rect -32 2730 4984 2740
rect -32 2690 40 2730
rect 4890 2690 4984 2730
rect -32 2674 4984 2690
rect -32 2660 34 2674
rect -32 790 -20 2660
rect 20 790 34 2660
rect 4918 2670 4984 2674
rect 1490 1170 4620 1200
rect 1490 1120 1530 1170
rect 4580 1120 4620 1170
rect 1490 1091 4620 1120
rect 1490 1090 1850 1091
rect 4260 1090 4620 1091
rect -32 760 34 790
rect 4918 780 4930 2670
rect 4970 780 4984 2670
rect 4918 760 4984 780
rect -32 750 4984 760
rect -32 710 40 750
rect 4900 710 4984 750
rect -32 694 4984 710
rect 6763 3015 7541 3049
rect 6763 2953 6797 3015
rect 5536 2834 5632 2868
rect 5770 2834 5866 2868
rect 5536 2772 5570 2834
rect 3496 72 3592 106
rect 5292 72 5388 106
rect 3496 10 3530 72
rect 5354 10 5388 72
rect 3496 -190 3530 -128
rect 5354 -190 5388 -128
rect 3496 -224 3592 -190
rect 5292 -224 5388 -190
rect 5832 2772 5866 2834
rect 5536 -190 5570 -128
rect 7507 2953 7541 3015
rect 6763 2597 6797 2659
rect 7507 2597 7541 2659
rect 6763 2563 6859 2597
rect 7445 2563 7541 2597
rect 6763 1555 7541 1589
rect 6763 1493 6797 1555
rect 7507 1493 7541 1555
rect 6763 1137 6797 1199
rect 7507 1137 7541 1199
rect 6763 1103 6859 1137
rect 7445 1103 7541 1137
rect 7415 173 7541 197
rect 7449 139 7507 173
rect 7415 92 7541 139
rect 5832 -190 5866 -128
rect 5536 -224 5632 -190
rect 5770 -224 5866 -190
<< nsubdiff >>
rect 6763 3583 6859 3617
rect 7445 3583 7541 3617
rect 6763 3520 6797 3583
rect 7507 3520 7541 3583
rect 6763 3155 6797 3218
rect 7507 3155 7541 3218
rect 6763 3121 7541 3155
rect -296 3060 5248 3070
rect -296 3020 -230 3060
rect 5170 3020 5248 3060
rect -296 3004 5248 3020
rect -296 2980 -230 3004
rect -296 450 -280 2980
rect -240 450 -230 2980
rect 5182 2990 5248 3004
rect 1530 2360 4620 2400
rect 1530 2320 1570 2360
rect 4580 2320 4620 2360
rect 1530 2290 4620 2320
rect -296 430 -230 450
rect 5182 440 5200 2990
rect 5240 440 5248 2990
rect 5182 430 5248 440
rect -296 420 5248 430
rect -296 380 -200 420
rect 5170 380 5248 420
rect -296 364 5248 380
rect 6763 2123 6859 2157
rect 7445 2123 7541 2157
rect 6763 2060 6797 2123
rect 7507 2060 7541 2123
rect 6763 1695 6797 1758
rect 7507 1695 7541 1758
rect 6763 1661 7541 1695
rect 7415 475 7541 508
rect 7449 441 7507 475
rect 7415 391 7541 441
rect 7449 357 7507 391
rect 7415 333 7541 357
<< psubdiffcont >>
rect 40 2690 4890 2730
rect -20 790 20 2660
rect 1530 1120 4580 1170
rect 4930 780 4970 2670
rect 40 710 4900 750
rect 5632 2834 5770 2868
rect 3592 72 5292 106
rect 3496 -128 3530 10
rect 5354 -128 5388 10
rect 3592 -224 5292 -190
rect 5536 -128 5570 2772
rect 5832 -128 5866 2772
rect 6763 2659 6797 2953
rect 7507 2659 7541 2953
rect 6859 2563 7445 2597
rect 6763 1199 6797 1493
rect 7507 1199 7541 1493
rect 6859 1103 7445 1137
rect 7415 139 7449 173
rect 7507 139 7541 173
rect 5632 -224 5770 -190
<< nsubdiffcont >>
rect 6859 3583 7445 3617
rect 6763 3218 6797 3520
rect 7507 3218 7541 3520
rect -230 3020 5170 3060
rect -280 450 -240 2980
rect 1570 2320 4580 2360
rect 5200 440 5240 2990
rect -200 380 5170 420
rect 6859 2123 7445 2157
rect 6763 1758 6797 2060
rect 7507 1758 7541 2060
rect 7415 441 7449 475
rect 7507 441 7541 475
rect 7415 357 7449 391
rect 7507 357 7541 391
<< poly >>
rect 6923 3514 7123 3530
rect 6923 3480 6939 3514
rect 7107 3480 7123 3514
rect 6923 3433 7123 3480
rect 7181 3514 7381 3530
rect 7181 3480 7197 3514
rect 7365 3480 7381 3514
rect 7181 3433 7381 3480
rect 6923 3207 7123 3233
rect 7181 3207 7381 3233
rect 1540 2232 1740 2258
rect 1798 2232 1998 2258
rect 2056 2232 2256 2258
rect 2314 2232 2514 2258
rect 2572 2232 2772 2258
rect 2830 2232 3030 2258
rect 3088 2232 3288 2258
rect 3346 2232 3546 2258
rect 3604 2232 3804 2258
rect 3862 2232 4062 2258
rect 4120 2232 4320 2258
rect 4378 2232 4578 2258
rect 1540 1985 1740 2032
rect 1540 1951 1556 1985
rect 1724 1951 1740 1985
rect 1540 1935 1740 1951
rect 1798 1985 1998 2032
rect 1798 1951 1814 1985
rect 1982 1951 1998 1985
rect 1798 1935 1998 1951
rect 2056 1985 2256 2032
rect 2056 1951 2072 1985
rect 2240 1951 2256 1985
rect 2056 1935 2256 1951
rect 2314 1985 2514 2032
rect 2314 1951 2330 1985
rect 2498 1951 2514 1985
rect 2314 1935 2514 1951
rect 2572 1985 2772 2032
rect 2572 1951 2588 1985
rect 2756 1951 2772 1985
rect 2572 1935 2772 1951
rect 2830 1985 3030 2032
rect 2830 1951 2846 1985
rect 3014 1951 3030 1985
rect 2830 1935 3030 1951
rect 3088 1985 3288 2032
rect 3088 1951 3104 1985
rect 3272 1951 3288 1985
rect 3088 1935 3288 1951
rect 3346 1985 3546 2032
rect 3346 1951 3362 1985
rect 3530 1951 3546 1985
rect 3346 1935 3546 1951
rect 3604 1985 3804 2032
rect 3604 1951 3620 1985
rect 3788 1951 3804 1985
rect 3604 1935 3804 1951
rect 3862 1985 4062 2032
rect 3862 1951 3878 1985
rect 4046 1951 4062 1985
rect 3862 1935 4062 1951
rect 4120 1985 4320 2032
rect 4120 1951 4136 1985
rect 4304 1951 4320 1985
rect 4120 1935 4320 1951
rect 4378 1985 4578 2032
rect 4378 1951 4394 1985
rect 4562 1951 4578 1985
rect 4378 1935 4578 1951
rect 1798 1877 1998 1893
rect 1798 1843 1814 1877
rect 1982 1843 1998 1877
rect 1540 1805 1740 1831
rect 1798 1805 1998 1843
rect 2572 1877 2772 1893
rect 2572 1843 2588 1877
rect 2756 1843 2772 1877
rect 2056 1805 2256 1831
rect 2314 1805 2514 1831
rect 2572 1805 2772 1843
rect 2830 1877 3030 1893
rect 2830 1843 2846 1877
rect 3014 1843 3030 1877
rect 2830 1805 3030 1843
rect 3604 1877 3804 1893
rect 3604 1843 3620 1877
rect 3788 1843 3804 1877
rect 3088 1805 3288 1831
rect 3346 1805 3546 1831
rect 3604 1805 3804 1843
rect 3862 1877 4062 1893
rect 3862 1843 3878 1877
rect 4046 1843 4062 1877
rect 3862 1805 4062 1843
rect 4120 1805 4320 1831
rect 4378 1805 4578 1831
rect 1540 1567 1740 1605
rect 1798 1579 1998 1605
rect 1540 1533 1556 1567
rect 1724 1533 1740 1567
rect 1540 1517 1740 1533
rect 2056 1567 2256 1605
rect 2056 1533 2072 1567
rect 2240 1533 2256 1567
rect 2056 1517 2256 1533
rect 2314 1567 2514 1605
rect 2572 1579 2772 1605
rect 2830 1579 3030 1605
rect 2314 1533 2330 1567
rect 2498 1533 2514 1567
rect 2314 1517 2514 1533
rect 3088 1567 3288 1605
rect 3088 1533 3104 1567
rect 3272 1533 3288 1567
rect 3088 1517 3288 1533
rect 3346 1567 3546 1605
rect 3604 1579 3804 1605
rect 3862 1579 4062 1605
rect 3346 1533 3362 1567
rect 3530 1533 3546 1567
rect 3346 1517 3546 1533
rect 4120 1567 4320 1605
rect 4120 1533 4136 1567
rect 4304 1533 4320 1567
rect 4120 1517 4320 1533
rect 4378 1567 4578 1605
rect 4378 1533 4394 1567
rect 4562 1533 4578 1567
rect 4378 1517 4578 1533
rect 1540 1441 1740 1457
rect 1540 1407 1556 1441
rect 1724 1407 1740 1441
rect 1540 1369 1740 1407
rect 1798 1441 1998 1457
rect 1798 1407 1814 1441
rect 1982 1407 1998 1441
rect 1798 1369 1998 1407
rect 2056 1441 2256 1457
rect 2056 1407 2072 1441
rect 2240 1407 2256 1441
rect 2056 1369 2256 1407
rect 2314 1441 2514 1457
rect 2314 1407 2330 1441
rect 2498 1407 2514 1441
rect 2314 1369 2514 1407
rect 2572 1441 2772 1457
rect 2572 1407 2588 1441
rect 2756 1407 2772 1441
rect 2572 1369 2772 1407
rect 2830 1441 3030 1457
rect 2830 1407 2846 1441
rect 3014 1407 3030 1441
rect 2830 1369 3030 1407
rect 3088 1441 3288 1457
rect 3088 1407 3104 1441
rect 3272 1407 3288 1441
rect 3088 1369 3288 1407
rect 3346 1441 3546 1457
rect 3346 1407 3362 1441
rect 3530 1407 3546 1441
rect 3346 1369 3546 1407
rect 3604 1441 3804 1457
rect 3604 1407 3620 1441
rect 3788 1407 3804 1441
rect 3604 1369 3804 1407
rect 3862 1441 4062 1457
rect 3862 1407 3878 1441
rect 4046 1407 4062 1441
rect 3862 1369 4062 1407
rect 4120 1441 4320 1457
rect 4120 1407 4136 1441
rect 4304 1407 4320 1441
rect 4120 1369 4320 1407
rect 4378 1441 4578 1457
rect 4378 1407 4394 1441
rect 4562 1407 4578 1441
rect 4378 1369 4578 1407
rect 1540 1259 1740 1285
rect 1798 1259 1998 1285
rect 2056 1259 2256 1285
rect 2314 1259 2514 1285
rect 2572 1259 2772 1285
rect 2830 1259 3030 1285
rect 3088 1259 3288 1285
rect 3346 1259 3546 1285
rect 3604 1259 3804 1285
rect 3862 1259 4062 1285
rect 4120 1259 4320 1285
rect 4378 1259 4578 1285
rect 6923 2937 7123 2963
rect 7181 2937 7381 2963
rect 6923 2699 7123 2737
rect 6923 2665 6939 2699
rect 7107 2665 7123 2699
rect 6923 2649 7123 2665
rect 7181 2699 7381 2737
rect 7181 2665 7197 2699
rect 7365 2665 7381 2699
rect 7181 2649 7381 2665
rect 6923 2054 7123 2070
rect 6923 2020 6939 2054
rect 7107 2020 7123 2054
rect 6923 1973 7123 2020
rect 7181 2054 7381 2070
rect 7181 2020 7197 2054
rect 7365 2020 7381 2054
rect 7181 1973 7381 2020
rect 6923 1747 7123 1773
rect 7181 1747 7381 1773
rect 6923 1477 7123 1503
rect 7181 1477 7381 1503
rect 6923 1239 7123 1277
rect 6923 1205 6939 1239
rect 7107 1205 7123 1239
rect 6923 1189 7123 1205
rect 7181 1239 7381 1277
rect 7181 1205 7197 1239
rect 7365 1205 7381 1239
rect 7181 1189 7381 1205
rect 6670 525 6700 551
rect 6754 525 6784 551
rect 6838 525 6868 551
rect 6922 525 6952 551
rect 7006 525 7036 551
rect 7090 525 7120 551
rect 7174 525 7204 551
rect 7258 525 7288 551
rect 6670 293 6700 325
rect 6754 293 6784 325
rect 6838 293 6868 325
rect 6922 293 6952 325
rect 7006 293 7036 325
rect 7090 293 7120 325
rect 7174 293 7204 325
rect 7258 293 7288 325
rect 6670 277 7288 293
rect 6670 243 6710 277
rect 6744 243 6794 277
rect 6828 243 6878 277
rect 6912 243 6962 277
rect 6996 243 7046 277
rect 7080 243 7130 277
rect 7164 243 7214 277
rect 7248 243 7288 277
rect 6670 227 7288 243
rect 6670 205 6700 227
rect 6754 205 6784 227
rect 6838 205 6868 227
rect 6922 205 6952 227
rect 7006 205 7036 227
rect 7090 205 7120 227
rect 7174 205 7204 227
rect 7258 205 7288 227
rect 6670 49 6700 75
rect 6754 49 6784 75
rect 6838 49 6868 75
rect 6922 49 6952 75
rect 7006 49 7036 75
rect 7090 49 7120 75
rect 7174 49 7204 75
rect 7258 49 7288 75
<< polycont >>
rect 6939 3480 7107 3514
rect 7197 3480 7365 3514
rect 1556 1951 1724 1985
rect 1814 1951 1982 1985
rect 2072 1951 2240 1985
rect 2330 1951 2498 1985
rect 2588 1951 2756 1985
rect 2846 1951 3014 1985
rect 3104 1951 3272 1985
rect 3362 1951 3530 1985
rect 3620 1951 3788 1985
rect 3878 1951 4046 1985
rect 4136 1951 4304 1985
rect 4394 1951 4562 1985
rect 1814 1843 1982 1877
rect 2588 1843 2756 1877
rect 2846 1843 3014 1877
rect 3620 1843 3788 1877
rect 3878 1843 4046 1877
rect 1556 1533 1724 1567
rect 2072 1533 2240 1567
rect 2330 1533 2498 1567
rect 3104 1533 3272 1567
rect 3362 1533 3530 1567
rect 4136 1533 4304 1567
rect 4394 1533 4562 1567
rect 1556 1407 1724 1441
rect 1814 1407 1982 1441
rect 2072 1407 2240 1441
rect 2330 1407 2498 1441
rect 2588 1407 2756 1441
rect 2846 1407 3014 1441
rect 3104 1407 3272 1441
rect 3362 1407 3530 1441
rect 3620 1407 3788 1441
rect 3878 1407 4046 1441
rect 4136 1407 4304 1441
rect 4394 1407 4562 1441
rect 6939 2665 7107 2699
rect 7197 2665 7365 2699
rect 6939 2020 7107 2054
rect 7197 2020 7365 2054
rect 6939 1205 7107 1239
rect 7197 1205 7365 1239
rect 6710 243 6744 277
rect 6794 243 6828 277
rect 6878 243 6912 277
rect 6962 243 6996 277
rect 7046 243 7080 277
rect 7130 243 7164 277
rect 7214 243 7248 277
<< xpolycontact >>
rect 896 2312 1328 2382
rect 896 1150 1328 1220
rect 3626 -94 4058 -24
rect 4826 -94 5258 -24
rect 5666 2306 5736 2738
rect 5666 -94 5736 338
<< xpolyres >>
rect 192 2312 896 2382
rect 192 2216 262 2312
rect 192 2146 792 2216
rect 722 2050 792 2146
rect 192 1980 792 2050
rect 192 1884 262 1980
rect 192 1814 792 1884
rect 722 1718 792 1814
rect 192 1648 792 1718
rect 192 1552 262 1648
rect 192 1482 792 1552
rect 722 1386 792 1482
rect 192 1316 792 1386
rect 192 1220 262 1316
rect 192 1150 896 1220
rect 4058 -94 4826 -24
rect 5666 338 5736 2306
<< locali >>
rect 6730 3617 7580 3630
rect 6730 3583 6859 3617
rect 7445 3583 7580 3617
rect 6730 3580 7580 3583
rect 6730 3520 6800 3580
rect 6730 3218 6763 3520
rect 6797 3218 6800 3520
rect 7500 3520 7580 3580
rect 6923 3480 6939 3514
rect 7107 3480 7123 3514
rect 7181 3480 7197 3514
rect 7365 3480 7381 3514
rect 6877 3430 6911 3437
rect 6730 3180 6800 3218
rect 6860 3421 6930 3430
rect 6860 3245 6877 3421
rect 6911 3260 6930 3421
rect 7135 3421 7169 3437
rect 7393 3430 7427 3437
rect 6911 3245 7060 3260
rect 6860 3180 7060 3245
rect 7380 3421 7440 3430
rect 7380 3260 7393 3421
rect 7135 3229 7169 3245
rect 7240 3245 7393 3260
rect 7427 3245 7440 3421
rect 7000 3100 7060 3180
rect 7240 3180 7440 3245
rect 7500 3218 7507 3520
rect 7541 3460 7580 3520
rect 7541 3420 7780 3460
rect 7541 3240 7660 3420
rect 7760 3240 7780 3420
rect 7541 3218 7780 3240
rect 7500 3200 7780 3218
rect 7240 3100 7300 3180
rect -296 3060 5248 3070
rect -296 380 -280 3060
rect -240 3004 5200 3020
rect -240 430 -230 3004
rect -32 2730 4984 2740
rect -32 710 -20 2730
rect 20 2674 4930 2690
rect 20 760 34 2674
rect 894 2382 4630 2400
rect 894 2312 896 2382
rect 1328 2360 4630 2382
rect 4580 2320 4630 2360
rect 1328 2312 4630 2320
rect 894 2280 4630 2312
rect 1494 2220 1528 2236
rect 1494 2028 1528 2044
rect 1752 2220 1786 2236
rect 1752 2028 1786 2044
rect 2010 2220 2044 2236
rect 2010 2028 2044 2044
rect 2268 2220 2302 2236
rect 2268 2028 2302 2044
rect 2526 2220 2560 2236
rect 2526 2028 2560 2044
rect 2784 2220 2818 2236
rect 2784 2028 2818 2044
rect 3042 2220 3076 2236
rect 3042 2028 3076 2044
rect 3300 2220 3334 2236
rect 3300 2028 3334 2044
rect 3558 2220 3592 2236
rect 3558 2028 3592 2044
rect 3816 2220 3850 2236
rect 3816 2028 3850 2044
rect 4074 2220 4108 2236
rect 4074 2028 4108 2044
rect 4332 2220 4366 2236
rect 4332 2028 4366 2044
rect 4590 2220 4624 2236
rect 4590 2028 4624 2044
rect 1540 1951 1556 1985
rect 1724 1951 1740 1985
rect 1798 1951 1814 1985
rect 1982 1951 1998 1985
rect 2056 1951 2072 1985
rect 2240 1951 2256 1985
rect 2314 1951 2330 1985
rect 2498 1951 2514 1985
rect 2572 1951 2588 1985
rect 2756 1951 2772 1985
rect 2830 1951 2846 1985
rect 3014 1951 3030 1985
rect 3088 1951 3104 1985
rect 3272 1951 3288 1985
rect 3346 1951 3362 1985
rect 3530 1951 3546 1985
rect 3604 1951 3620 1985
rect 3788 1951 3804 1985
rect 3862 1951 3878 1985
rect 4046 1951 4062 1985
rect 4120 1951 4136 1985
rect 4304 1951 4320 1985
rect 4378 1951 4394 1985
rect 4562 1951 4578 1985
rect 1798 1843 1814 1877
rect 1982 1843 1998 1877
rect 2572 1843 2588 1877
rect 2756 1843 2772 1877
rect 2830 1843 2846 1877
rect 3014 1843 3030 1877
rect 3604 1843 3620 1877
rect 3788 1843 3804 1877
rect 3862 1843 3878 1877
rect 4046 1843 4062 1877
rect 1494 1793 1528 1809
rect 1494 1601 1528 1617
rect 1752 1793 1786 1809
rect 1752 1601 1786 1617
rect 2010 1793 2044 1809
rect 2010 1601 2044 1617
rect 2268 1793 2302 1809
rect 2268 1601 2302 1617
rect 2526 1793 2560 1809
rect 2526 1601 2560 1617
rect 2784 1793 2818 1809
rect 2784 1601 2818 1617
rect 3042 1793 3076 1809
rect 3042 1601 3076 1617
rect 3300 1793 3334 1809
rect 3300 1601 3334 1617
rect 3558 1793 3592 1809
rect 3558 1601 3592 1617
rect 3816 1793 3850 1809
rect 3816 1601 3850 1617
rect 4074 1793 4108 1809
rect 4074 1601 4108 1617
rect 4332 1793 4366 1809
rect 4332 1601 4366 1617
rect 4590 1793 4624 1809
rect 4590 1601 4624 1617
rect 1540 1533 1556 1567
rect 1724 1533 1740 1567
rect 2056 1533 2072 1567
rect 2240 1533 2256 1567
rect 2314 1533 2330 1567
rect 2498 1533 2514 1567
rect 3088 1533 3104 1567
rect 3272 1533 3288 1567
rect 3346 1533 3362 1567
rect 3530 1533 3546 1567
rect 4120 1533 4136 1567
rect 4304 1533 4320 1567
rect 4378 1533 4394 1567
rect 4562 1533 4578 1567
rect 1540 1407 1556 1441
rect 1724 1407 1740 1441
rect 1798 1407 1814 1441
rect 1982 1407 1998 1441
rect 2056 1407 2072 1441
rect 2240 1407 2256 1441
rect 2314 1407 2330 1441
rect 2498 1407 2514 1441
rect 2572 1407 2588 1441
rect 2756 1407 2772 1441
rect 2830 1407 2846 1441
rect 3014 1407 3030 1441
rect 3088 1407 3104 1441
rect 3272 1407 3288 1441
rect 3346 1407 3362 1441
rect 3530 1407 3546 1441
rect 3604 1407 3620 1441
rect 3788 1407 3804 1441
rect 3862 1407 3878 1441
rect 4046 1407 4062 1441
rect 4120 1407 4136 1441
rect 4304 1407 4320 1441
rect 4378 1407 4394 1441
rect 4562 1407 4578 1441
rect 1494 1357 1528 1373
rect 1494 1281 1528 1297
rect 1752 1357 1786 1373
rect 1752 1281 1786 1297
rect 2010 1357 2044 1373
rect 2010 1281 2044 1297
rect 2268 1357 2302 1373
rect 2268 1281 2302 1297
rect 2526 1357 2560 1373
rect 2526 1281 2560 1297
rect 2784 1357 2818 1373
rect 2784 1281 2818 1297
rect 3042 1357 3076 1373
rect 3042 1281 3076 1297
rect 3300 1357 3334 1373
rect 3300 1281 3334 1297
rect 3558 1357 3592 1373
rect 3558 1281 3592 1297
rect 3816 1357 3850 1373
rect 3816 1281 3850 1297
rect 4074 1357 4108 1373
rect 4074 1281 4108 1297
rect 4332 1357 4366 1373
rect 4332 1281 4366 1297
rect 4590 1357 4624 1373
rect 4590 1281 4624 1297
rect 894 1230 1380 1260
rect 894 1220 960 1230
rect 894 1150 896 1220
rect 894 1140 960 1150
rect 1360 1140 1380 1230
rect 894 1120 1380 1140
rect 1490 1170 4630 1200
rect 1490 1120 1530 1170
rect 4580 1120 4630 1170
rect 1490 1090 4630 1120
rect 4918 760 4930 2674
rect 20 750 4930 760
rect 4970 710 4984 2730
rect -32 694 4984 710
rect 5182 430 5200 3004
rect -240 420 5200 430
rect 5240 380 5248 3060
rect 7000 3020 7300 3100
rect 6730 2953 6800 2980
rect 5536 2834 5632 2868
rect 5770 2834 5866 2868
rect 5536 2772 5570 2834
rect 5420 1180 5536 1200
rect 5832 2772 5866 2834
rect 5620 2738 5780 2740
rect 5620 2720 5666 2738
rect 5736 2720 5780 2738
rect 5620 2320 5640 2720
rect 5760 2320 5780 2720
rect 5620 2306 5666 2320
rect 5736 2306 5780 2320
rect 5620 2300 5780 2306
rect 5420 740 5440 1180
rect 5420 720 5536 740
rect -296 364 5248 380
rect 3520 180 4680 200
rect 3520 106 3540 180
rect 4660 106 4680 180
rect 3496 100 3540 106
rect 5292 100 5388 106
rect 3496 72 3592 100
rect 5292 72 5536 100
rect 3496 10 3530 72
rect 5354 10 5536 72
rect 3496 -190 3530 -128
rect 5388 -128 5536 10
rect 5354 -190 5570 -128
rect 6730 2659 6763 2953
rect 6797 2659 6800 2953
rect 6860 2925 6930 2980
rect 6860 2780 6877 2925
rect 6911 2780 6930 2925
rect 7100 2925 7200 3020
rect 6877 2733 6911 2749
rect 7100 2749 7135 2925
rect 7169 2749 7200 2925
rect 7380 2925 7440 2980
rect 7380 2780 7393 2925
rect 7100 2740 7200 2749
rect 7427 2780 7440 2925
rect 7500 2953 7780 2980
rect 7135 2733 7169 2740
rect 7393 2733 7427 2749
rect 6923 2665 6939 2699
rect 7107 2665 7123 2699
rect 7181 2665 7197 2699
rect 7365 2665 7381 2699
rect 6730 2600 6800 2659
rect 7500 2659 7507 2953
rect 7541 2940 7780 2953
rect 7541 2760 7660 2940
rect 7760 2760 7780 2940
rect 7541 2720 7780 2760
rect 7541 2659 7580 2720
rect 7500 2600 7580 2659
rect 6730 2597 7580 2600
rect 6730 2563 6859 2597
rect 7445 2563 7580 2597
rect 6730 2530 7580 2563
rect 6730 2157 7580 2170
rect 6730 2123 6859 2157
rect 7445 2123 7580 2157
rect 6730 2120 7580 2123
rect 6730 2060 6800 2120
rect 6730 1758 6763 2060
rect 6797 1758 6800 2060
rect 7500 2060 7580 2120
rect 6923 2020 6939 2054
rect 7107 2020 7123 2054
rect 7181 2020 7197 2054
rect 7365 2020 7381 2054
rect 6877 1970 6911 1977
rect 6730 1720 6800 1758
rect 6860 1961 6930 1970
rect 6860 1785 6877 1961
rect 6911 1800 6930 1961
rect 7135 1961 7169 1977
rect 7393 1970 7427 1977
rect 6911 1785 7060 1800
rect 6860 1720 7060 1785
rect 7380 1961 7440 1970
rect 7380 1800 7393 1961
rect 7135 1769 7169 1785
rect 7240 1785 7393 1800
rect 7427 1785 7440 1961
rect 7000 1640 7060 1720
rect 7240 1720 7440 1785
rect 7500 1758 7507 2060
rect 7541 2000 7580 2060
rect 7541 1960 7780 2000
rect 7541 1780 7660 1960
rect 7760 1780 7780 1960
rect 7541 1758 7780 1780
rect 7500 1740 7780 1758
rect 7240 1640 7300 1720
rect 7000 1560 7300 1640
rect 6730 1493 6800 1520
rect 6730 1199 6763 1493
rect 6797 1199 6800 1493
rect 6860 1465 6930 1520
rect 6860 1320 6877 1465
rect 6911 1320 6930 1465
rect 7100 1465 7200 1560
rect 6877 1273 6911 1289
rect 7100 1289 7135 1465
rect 7169 1289 7200 1465
rect 7380 1465 7440 1520
rect 7380 1320 7393 1465
rect 7100 1280 7200 1289
rect 7427 1320 7440 1465
rect 7500 1493 7780 1520
rect 7135 1273 7169 1280
rect 7393 1273 7427 1289
rect 6923 1205 6939 1239
rect 7107 1205 7123 1239
rect 7181 1205 7197 1239
rect 7365 1205 7381 1239
rect 6730 1140 6800 1199
rect 7500 1199 7507 1493
rect 7541 1480 7780 1493
rect 7541 1300 7660 1480
rect 7760 1300 7780 1480
rect 7541 1260 7780 1300
rect 7541 1199 7580 1260
rect 7500 1140 7580 1199
rect 6730 1137 7580 1140
rect 6730 1103 6859 1137
rect 7445 1103 7580 1137
rect 6730 1070 7580 1103
rect 6558 555 6587 589
rect 6621 555 6679 589
rect 6713 555 6771 589
rect 6805 555 6863 589
rect 6897 555 6955 589
rect 6989 555 7047 589
rect 7081 555 7139 589
rect 7173 555 7231 589
rect 7265 555 7323 589
rect 7357 555 7415 589
rect 7449 555 7507 589
rect 7541 555 7570 589
rect 6609 513 6660 555
rect 6609 479 6626 513
rect 6609 445 6660 479
rect 6609 411 6626 445
rect 6609 395 6660 411
rect 6694 513 6760 521
rect 6694 479 6710 513
rect 6744 479 6760 513
rect 6694 445 6760 479
rect 6694 411 6710 445
rect 6744 411 6760 445
rect 6694 377 6760 411
rect 6794 513 6828 555
rect 6794 445 6828 479
rect 6794 395 6828 411
rect 6862 513 6928 521
rect 6862 479 6878 513
rect 6912 479 6928 513
rect 6862 445 6928 479
rect 6862 411 6878 445
rect 6912 411 6928 445
rect 6694 361 6710 377
rect 6575 343 6710 361
rect 6744 361 6760 377
rect 6862 377 6928 411
rect 6962 513 6996 555
rect 6962 445 6996 479
rect 6962 395 6996 411
rect 7030 513 7096 521
rect 7030 479 7046 513
rect 7080 479 7096 513
rect 7030 445 7096 479
rect 7030 411 7046 445
rect 7080 411 7096 445
rect 6862 361 6878 377
rect 6744 343 6878 361
rect 6912 361 6928 377
rect 7030 377 7096 411
rect 7130 513 7164 555
rect 7130 445 7164 479
rect 7130 395 7164 411
rect 7198 513 7264 521
rect 7198 479 7214 513
rect 7248 479 7264 513
rect 7198 445 7264 479
rect 7198 411 7214 445
rect 7248 411 7264 445
rect 7030 361 7046 377
rect 6912 343 7046 361
rect 7080 361 7096 377
rect 7198 377 7264 411
rect 7298 513 7358 555
rect 7332 479 7358 513
rect 7298 445 7358 479
rect 7332 411 7358 445
rect 7298 395 7358 411
rect 7403 475 7553 519
rect 7403 441 7415 475
rect 7449 441 7507 475
rect 7541 441 7553 475
rect 7198 361 7214 377
rect 7080 343 7214 361
rect 7248 361 7264 377
rect 7403 391 7553 441
rect 7248 348 7369 361
rect 7248 343 7314 348
rect 6575 327 7314 343
rect 6575 209 6644 327
rect 6694 284 7265 293
rect 6694 250 6702 284
rect 7190 277 7265 284
rect 7190 250 7214 277
rect 6694 243 6710 250
rect 6744 243 6794 250
rect 6828 243 6878 250
rect 6912 243 6962 250
rect 6996 243 7046 250
rect 7080 243 7130 250
rect 7164 243 7214 250
rect 7248 243 7265 277
rect 7305 209 7314 327
rect 6575 189 7314 209
rect 6575 171 6710 189
rect 6694 155 6710 171
rect 6744 171 6878 189
rect 6744 155 6760 171
rect 6609 121 6660 137
rect 6609 87 6626 121
rect 6609 45 6660 87
rect 6694 121 6760 155
rect 6862 155 6878 171
rect 6912 171 7046 189
rect 6912 155 6928 171
rect 6694 87 6710 121
rect 6744 87 6760 121
rect 6694 79 6760 87
rect 6794 121 6828 137
rect 6794 45 6828 87
rect 6862 121 6928 155
rect 7030 155 7046 171
rect 7080 171 7214 189
rect 7080 155 7096 171
rect 6862 87 6878 121
rect 6912 87 6928 121
rect 6862 79 6928 87
rect 6962 121 6996 137
rect 6962 45 6996 87
rect 7030 121 7096 155
rect 7198 155 7214 171
rect 7248 184 7314 189
rect 7362 184 7369 348
rect 7403 357 7415 391
rect 7449 357 7507 391
rect 7541 357 7553 391
rect 7403 322 7553 357
rect 7248 171 7369 184
rect 7403 173 7553 190
rect 7248 155 7264 171
rect 7030 87 7046 121
rect 7080 87 7096 121
rect 7030 79 7096 87
rect 7130 121 7164 137
rect 7130 45 7164 87
rect 7198 121 7264 155
rect 7403 139 7415 173
rect 7449 139 7507 173
rect 7541 139 7553 173
rect 7198 87 7214 121
rect 7248 87 7264 121
rect 7198 79 7264 87
rect 7298 121 7359 137
rect 7332 87 7359 121
rect 7298 45 7359 87
rect 7403 81 7553 139
rect 6558 11 6587 45
rect 6621 11 6679 45
rect 6713 11 6771 45
rect 6805 11 6863 45
rect 6897 11 6955 45
rect 6989 11 7047 45
rect 7081 11 7139 45
rect 7173 11 7231 45
rect 7265 11 7323 45
rect 7357 11 7415 45
rect 7449 11 7507 45
rect 7541 11 7570 45
rect 5832 -190 5866 -128
rect 3496 -224 3592 -190
rect 5292 -220 5632 -190
rect 5292 -224 5388 -220
rect 5536 -224 5632 -220
rect 5770 -224 5866 -190
<< viali >>
rect 6939 3480 7107 3514
rect 7197 3480 7365 3514
rect 6877 3245 6911 3421
rect 7135 3245 7169 3421
rect 7393 3245 7427 3421
rect 7660 3240 7760 3420
rect -280 3020 -230 3060
rect -230 3020 5170 3060
rect 5170 3020 5240 3060
rect -280 2980 -240 3020
rect -280 450 -240 2980
rect -280 420 -240 450
rect -20 2690 40 2730
rect 40 2690 4890 2730
rect 4890 2690 4970 2730
rect -20 2660 20 2690
rect -20 790 20 2660
rect -20 750 20 790
rect 1000 2320 1328 2360
rect 1328 2320 1570 2360
rect 1570 2320 4580 2360
rect 1494 2044 1528 2220
rect 1752 2044 1786 2220
rect 2010 2044 2044 2220
rect 2268 2044 2302 2220
rect 2526 2044 2560 2220
rect 2784 2044 2818 2220
rect 3042 2044 3076 2220
rect 3300 2044 3334 2220
rect 3558 2044 3592 2220
rect 3816 2044 3850 2220
rect 4074 2044 4108 2220
rect 4332 2044 4366 2220
rect 4590 2044 4624 2220
rect 1556 1951 1724 1985
rect 1814 1951 1982 1985
rect 2072 1951 2240 1985
rect 2330 1951 2498 1985
rect 2588 1951 2756 1985
rect 2846 1951 3014 1985
rect 3104 1951 3272 1985
rect 3362 1951 3530 1985
rect 3620 1951 3788 1985
rect 3878 1951 4046 1985
rect 4136 1951 4304 1985
rect 4394 1951 4562 1985
rect 1814 1843 1982 1877
rect 2588 1843 2756 1877
rect 2846 1843 3014 1877
rect 3620 1843 3788 1877
rect 3878 1843 4046 1877
rect 1494 1617 1528 1793
rect 1752 1617 1786 1793
rect 2010 1617 2044 1793
rect 2268 1617 2302 1793
rect 2526 1617 2560 1793
rect 2784 1617 2818 1793
rect 3042 1617 3076 1793
rect 3300 1617 3334 1793
rect 3558 1617 3592 1793
rect 3816 1617 3850 1793
rect 4074 1617 4108 1793
rect 4332 1617 4366 1793
rect 4590 1617 4624 1793
rect 1556 1533 1724 1567
rect 2072 1533 2240 1567
rect 2330 1533 2498 1567
rect 3104 1533 3272 1567
rect 3362 1533 3530 1567
rect 4136 1533 4304 1567
rect 4394 1533 4562 1567
rect 1556 1407 1724 1441
rect 1814 1407 1982 1441
rect 2072 1407 2240 1441
rect 2330 1407 2498 1441
rect 2588 1407 2756 1441
rect 2846 1407 3014 1441
rect 3104 1407 3272 1441
rect 3362 1407 3530 1441
rect 3620 1407 3788 1441
rect 3878 1407 4046 1441
rect 4136 1407 4304 1441
rect 4394 1407 4562 1441
rect 1494 1297 1528 1357
rect 1752 1297 1786 1357
rect 2010 1297 2044 1357
rect 2268 1297 2302 1357
rect 2526 1297 2560 1357
rect 2784 1297 2818 1357
rect 3042 1297 3076 1357
rect 3300 1297 3334 1357
rect 3558 1297 3592 1357
rect 3816 1297 3850 1357
rect 4074 1297 4108 1357
rect 4332 1297 4366 1357
rect 4590 1297 4624 1357
rect 960 1220 1360 1230
rect 960 1150 1328 1220
rect 1328 1150 1360 1220
rect 960 1140 1360 1150
rect 1530 1120 4580 1170
rect 4930 2670 4970 2690
rect 4930 780 4970 2670
rect 4930 750 4970 780
rect -20 710 40 750
rect 40 710 4900 750
rect 4900 710 4970 750
rect 5200 2990 5240 3020
rect 5200 440 5240 2990
rect 5200 420 5240 440
rect -280 380 -200 420
rect -200 380 5170 420
rect 5170 380 5240 420
rect 5640 2320 5666 2720
rect 5666 2320 5736 2720
rect 5736 2320 5760 2720
rect 5440 740 5536 1180
rect 5536 740 5540 1180
rect 3540 106 4660 180
rect 3540 100 3592 106
rect 3592 100 4660 106
rect 3644 -78 4041 -40
rect 4843 -78 5240 -40
rect 5682 -76 5720 321
rect 6877 2749 6911 2925
rect 7135 2749 7169 2925
rect 7393 2749 7427 2925
rect 6939 2665 7107 2699
rect 7197 2665 7365 2699
rect 7660 2760 7760 2940
rect 6939 2020 7107 2054
rect 7197 2020 7365 2054
rect 6877 1785 6911 1961
rect 7135 1785 7169 1961
rect 7393 1785 7427 1961
rect 7660 1780 7760 1960
rect 6877 1289 6911 1465
rect 7135 1289 7169 1465
rect 7393 1289 7427 1465
rect 6939 1205 7107 1239
rect 7197 1205 7365 1239
rect 7660 1300 7760 1480
rect 6587 555 6621 589
rect 6679 555 6713 589
rect 6771 555 6805 589
rect 6863 555 6897 589
rect 6955 555 6989 589
rect 7047 555 7081 589
rect 7139 555 7173 589
rect 7231 555 7265 589
rect 7323 555 7357 589
rect 7415 555 7449 589
rect 7507 555 7541 589
rect 6702 277 7190 284
rect 6702 250 6710 277
rect 6710 250 6744 277
rect 6744 250 6794 277
rect 6794 250 6828 277
rect 6828 250 6878 277
rect 6878 250 6912 277
rect 6912 250 6962 277
rect 6962 250 6996 277
rect 6996 250 7046 277
rect 7046 250 7080 277
rect 7080 250 7130 277
rect 7130 250 7164 277
rect 7164 250 7190 277
rect 7314 184 7362 348
rect 6587 11 6621 45
rect 6679 11 6713 45
rect 6771 11 6805 45
rect 6863 11 6897 45
rect 6955 11 6989 45
rect 7047 11 7081 45
rect 7139 11 7173 45
rect 7231 11 7265 45
rect 7323 11 7357 45
rect 7415 11 7449 45
rect 7507 11 7541 45
<< metal1 >>
rect 6920 3760 7380 3780
rect 6920 3580 6940 3760
rect 7360 3580 7380 3760
rect 6920 3514 7380 3580
rect 6920 3480 6939 3514
rect 7107 3480 7197 3514
rect 7365 3480 7380 3514
rect 6927 3474 7119 3480
rect 7185 3474 7377 3480
rect 7840 3440 8680 3480
rect 6700 3421 6960 3440
rect 6700 3420 6877 3421
rect 6911 3420 6960 3421
rect 6700 3240 6720 3420
rect 6940 3240 6960 3420
rect 6700 3220 6960 3240
rect 7100 3421 7200 3440
rect 7100 3245 7135 3421
rect 7169 3245 7200 3421
rect 7100 3140 7200 3245
rect 7340 3421 7600 3440
rect 7340 3420 7393 3421
rect 7427 3420 7600 3421
rect 7340 3240 7360 3420
rect 7580 3240 7600 3420
rect 7340 3220 7600 3240
rect 7640 3420 8680 3440
rect 7640 3240 7660 3420
rect 7760 3240 8560 3420
rect 7640 3220 8560 3240
rect 7840 3200 8560 3220
rect 8640 3200 8680 3420
rect 7840 3180 8680 3200
rect -380 3100 5320 3120
rect -380 3060 1450 3100
rect 4660 3060 5320 3100
rect -380 380 -280 3060
rect -240 2940 1450 3020
rect 4660 2940 5200 3020
rect -240 2920 5200 2940
rect -240 520 -180 2920
rect -80 2730 5020 2820
rect -80 710 -20 2730
rect 20 2620 4930 2690
rect 20 820 120 2620
rect 894 2380 4630 2400
rect 894 2360 1450 2380
rect 894 2320 1000 2360
rect 894 2300 1450 2320
rect 4610 2300 4630 2380
rect 894 2280 4630 2300
rect 1490 2232 1550 2280
rect 1488 2220 1550 2232
rect 1740 2230 1800 2240
rect 1488 2044 1494 2220
rect 1528 2044 1550 2220
rect 1488 2032 1550 2044
rect 1700 2220 1850 2230
rect 1700 2110 1752 2220
rect 1786 2110 1850 2220
rect 1700 2050 1710 2110
rect 1820 2050 1850 2110
rect 1700 2044 1752 2050
rect 1786 2044 1850 2050
rect 1700 2040 1850 2044
rect 1960 2220 2090 2280
rect 2262 2230 2308 2232
rect 1960 2044 2010 2220
rect 2044 2044 2090 2220
rect 1960 2040 2090 2044
rect 2220 2220 2350 2230
rect 2220 2110 2268 2220
rect 2302 2110 2350 2220
rect 2220 2050 2230 2110
rect 2340 2050 2350 2110
rect 2220 2044 2268 2050
rect 2302 2044 2350 2050
rect 2220 2040 2350 2044
rect 2480 2220 2610 2280
rect 2480 2044 2526 2220
rect 2560 2044 2610 2220
rect 2480 2040 2610 2044
rect 2730 2220 2860 2240
rect 2730 2110 2784 2220
rect 2818 2110 2860 2220
rect 1490 1991 1550 2032
rect 1740 2030 1850 2040
rect 2004 2032 2050 2040
rect 2262 2032 2308 2040
rect 2520 2032 2566 2040
rect 1800 1991 1850 2030
rect 2730 2000 2740 2110
rect 2850 2000 2860 2110
rect 2990 2220 3120 2280
rect 3294 2230 3340 2232
rect 2990 2044 3042 2220
rect 3076 2044 3120 2220
rect 2990 2040 3120 2044
rect 3250 2220 3380 2230
rect 3250 2120 3300 2220
rect 3334 2120 3380 2220
rect 3250 2050 3260 2120
rect 3370 2050 3380 2120
rect 3250 2044 3300 2050
rect 3334 2044 3380 2050
rect 3250 2040 3380 2044
rect 3510 2220 3640 2280
rect 3510 2044 3558 2220
rect 3592 2044 3640 2220
rect 3510 2040 3640 2044
rect 3770 2220 3900 2240
rect 3770 2120 3816 2220
rect 3850 2120 3900 2220
rect 3036 2032 3082 2040
rect 3294 2032 3340 2040
rect 3552 2032 3598 2040
rect 2730 1991 2860 2000
rect 3770 2000 3780 2120
rect 3890 2000 3900 2120
rect 4030 2220 4160 2280
rect 4590 2232 4630 2280
rect 4326 2230 4372 2232
rect 4030 2044 4074 2220
rect 4108 2044 4160 2220
rect 4030 2040 4160 2044
rect 4280 2220 4410 2230
rect 4280 2120 4332 2220
rect 4366 2120 4410 2220
rect 4280 2050 4290 2120
rect 4400 2050 4410 2120
rect 4280 2044 4332 2050
rect 4366 2044 4410 2050
rect 4280 2040 4410 2044
rect 4584 2220 4630 2232
rect 4584 2044 4590 2220
rect 4624 2044 4630 2220
rect 4068 2032 4114 2040
rect 4326 2032 4372 2040
rect 4584 2032 4630 2044
rect 4590 2000 4630 2032
rect 3770 1991 3900 2000
rect 1490 1990 1736 1991
rect 1490 1985 1740 1990
rect 1800 1985 1994 1991
rect 2060 1985 2252 1991
rect 2318 1985 2510 1991
rect 2576 1985 3026 1991
rect 3092 1985 3284 1991
rect 3350 1985 3542 1991
rect 3608 1985 4058 1991
rect 4124 1985 4316 1991
rect 4380 1985 4630 2000
rect 1490 1951 1556 1985
rect 1724 1951 1740 1985
rect 1798 1951 1814 1985
rect 1982 1951 2072 1985
rect 2240 1951 2330 1985
rect 2498 1951 2588 1985
rect 2756 1951 2846 1985
rect 3014 1951 3104 1985
rect 3272 1951 3362 1985
rect 3530 1951 3620 1985
rect 3788 1951 3878 1985
rect 4046 1951 4136 1985
rect 4304 1951 4320 1985
rect 4380 1951 4394 1985
rect 4562 1951 4630 1985
rect 1490 1950 1740 1951
rect 1800 1950 1994 1951
rect 1544 1945 1736 1950
rect 1802 1945 1994 1950
rect 2060 1945 2252 1951
rect 2318 1945 2510 1951
rect 2576 1945 2768 1951
rect 2834 1945 3026 1951
rect 3092 1945 3284 1951
rect 3350 1945 3542 1951
rect 3608 1945 3800 1951
rect 3866 1945 4058 1951
rect 4124 1945 4316 1951
rect 4380 1950 4630 1951
rect 4382 1945 4574 1950
rect 2080 1900 2190 1910
rect 1802 1877 1994 1883
rect 2080 1877 2090 1900
rect 1798 1843 1814 1877
rect 1982 1843 2090 1877
rect 1802 1837 1994 1843
rect 1490 1805 1540 1810
rect 1488 1793 1540 1805
rect 1746 1800 1792 1805
rect 1488 1617 1494 1793
rect 1528 1617 1540 1793
rect 1488 1605 1540 1617
rect 1700 1793 1830 1800
rect 1700 1790 1752 1793
rect 1786 1790 1830 1793
rect 1700 1730 1710 1790
rect 1820 1730 1830 1790
rect 1700 1617 1752 1730
rect 1786 1617 1830 1730
rect 2004 1793 2050 1805
rect 2004 1700 2010 1793
rect 1700 1610 1830 1617
rect 1960 1680 2010 1700
rect 2044 1700 2050 1793
rect 2080 1740 2090 1843
rect 2180 1877 2190 1900
rect 4150 1900 4250 1910
rect 2576 1877 2768 1883
rect 2834 1877 3026 1883
rect 3608 1877 3800 1883
rect 3866 1877 4058 1883
rect 2180 1843 2588 1877
rect 2756 1843 2846 1877
rect 3014 1843 3620 1877
rect 3788 1843 3878 1877
rect 4046 1843 4062 1877
rect 2180 1740 2190 1843
rect 2576 1837 2768 1843
rect 2834 1837 3026 1843
rect 3608 1837 3800 1843
rect 3866 1837 4058 1843
rect 2262 1800 2308 1805
rect 2520 1800 2566 1805
rect 2778 1800 2824 1805
rect 3036 1800 3082 1805
rect 3294 1800 3340 1805
rect 3552 1800 3598 1805
rect 3810 1800 3856 1805
rect 2080 1730 2190 1740
rect 2220 1793 2350 1800
rect 2220 1790 2268 1793
rect 2302 1790 2350 1793
rect 2220 1730 2230 1790
rect 2340 1730 2350 1790
rect 2044 1680 2090 1700
rect 1960 1620 1970 1680
rect 2080 1620 2090 1680
rect 1960 1617 2010 1620
rect 2044 1617 2090 1620
rect 1960 1610 2090 1617
rect 2220 1617 2268 1730
rect 2302 1617 2350 1730
rect 2220 1610 2350 1617
rect 2480 1793 2610 1800
rect 2480 1680 2526 1793
rect 2560 1680 2610 1793
rect 2480 1620 2490 1680
rect 2600 1620 2610 1680
rect 2480 1617 2526 1620
rect 2560 1617 2610 1620
rect 2480 1610 2610 1617
rect 2730 1793 2860 1800
rect 2730 1790 2784 1793
rect 2818 1790 2860 1793
rect 2730 1730 2740 1790
rect 2850 1730 2860 1790
rect 2730 1617 2784 1730
rect 2818 1617 2860 1730
rect 2730 1610 2860 1617
rect 3000 1793 3130 1800
rect 3000 1680 3042 1793
rect 3076 1680 3130 1793
rect 3000 1620 3010 1680
rect 3120 1620 3130 1680
rect 3000 1617 3042 1620
rect 3076 1617 3130 1620
rect 3000 1610 3130 1617
rect 3250 1793 3380 1800
rect 3250 1790 3300 1793
rect 3334 1790 3380 1793
rect 3250 1730 3260 1790
rect 3370 1730 3380 1790
rect 3250 1617 3300 1730
rect 3334 1617 3380 1730
rect 3250 1610 3380 1617
rect 3510 1793 3640 1800
rect 3510 1680 3558 1793
rect 3592 1680 3640 1793
rect 3510 1620 3520 1680
rect 3630 1620 3640 1680
rect 3510 1617 3558 1620
rect 3592 1617 3640 1620
rect 3510 1610 3640 1617
rect 3770 1793 3900 1800
rect 3770 1790 3816 1793
rect 3850 1790 3900 1793
rect 3770 1730 3780 1790
rect 3890 1730 3900 1790
rect 3770 1617 3816 1730
rect 3850 1617 3900 1730
rect 4068 1793 4114 1805
rect 4068 1690 4074 1793
rect 3770 1610 3900 1617
rect 4020 1680 4074 1690
rect 4108 1690 4114 1793
rect 4150 1750 4160 1900
rect 4240 1750 4250 1900
rect 4326 1800 4372 1805
rect 4150 1720 4250 1750
rect 4108 1680 4150 1690
rect 4020 1620 4030 1680
rect 4140 1620 4150 1680
rect 4020 1617 4074 1620
rect 4108 1617 4150 1620
rect 4020 1610 4150 1617
rect 1746 1605 1792 1610
rect 2004 1605 2050 1610
rect 2262 1605 2308 1610
rect 2520 1605 2566 1610
rect 2778 1605 2824 1610
rect 3036 1605 3082 1610
rect 3294 1605 3340 1610
rect 3552 1605 3598 1610
rect 3810 1605 3856 1610
rect 4068 1605 4114 1610
rect 1490 1600 1540 1605
rect 1490 1573 1560 1600
rect 4180 1573 4250 1720
rect 4280 1793 4410 1800
rect 4280 1790 4332 1793
rect 4366 1790 4410 1793
rect 4280 1730 4290 1790
rect 4400 1730 4410 1790
rect 4280 1617 4332 1730
rect 4366 1617 4410 1730
rect 4280 1610 4410 1617
rect 4580 1793 4630 1810
rect 4580 1617 4590 1793
rect 4624 1617 4630 1793
rect 4326 1605 4372 1610
rect 4580 1600 4630 1617
rect 4550 1573 4630 1600
rect 1490 1570 1736 1573
rect 1490 1567 1740 1570
rect 2060 1567 2252 1573
rect 2318 1567 2510 1573
rect 3092 1567 3284 1573
rect 3350 1567 3542 1573
rect 4124 1567 4316 1573
rect 4382 1570 4630 1573
rect 4370 1567 4630 1570
rect 1490 1533 1556 1567
rect 1724 1533 1740 1567
rect 2056 1533 2072 1567
rect 2240 1533 2330 1567
rect 2498 1533 3104 1567
rect 3272 1533 3362 1567
rect 3530 1533 4136 1567
rect 4304 1533 4320 1567
rect 4370 1533 4394 1567
rect 4562 1533 4630 1567
rect 1490 1470 1740 1533
rect 2060 1527 2252 1533
rect 2318 1527 2510 1533
rect 3092 1527 3284 1533
rect 3350 1527 3542 1533
rect 4124 1527 4316 1533
rect 1490 1441 2260 1470
rect 2940 1460 2950 1490
rect 1490 1407 1556 1441
rect 1724 1407 1814 1441
rect 1982 1407 2072 1441
rect 2240 1407 2260 1441
rect 1490 1390 2260 1407
rect 2310 1441 2950 1460
rect 3170 1460 3180 1490
rect 4370 1470 4630 1533
rect 3170 1441 3810 1460
rect 2310 1407 2330 1441
rect 2498 1407 2588 1441
rect 2756 1407 2846 1441
rect 3014 1407 3104 1430
rect 3272 1407 3362 1441
rect 3530 1407 3620 1441
rect 3788 1407 3810 1441
rect 2310 1400 3810 1407
rect 3860 1441 4630 1470
rect 3860 1407 3878 1441
rect 4046 1407 4136 1441
rect 4304 1407 4394 1441
rect 4562 1407 4630 1441
rect 2940 1390 3180 1400
rect 1490 1370 2280 1390
rect 1490 1369 2304 1370
rect 1488 1357 2308 1369
rect 1488 1297 1494 1357
rect 1528 1297 1752 1357
rect 1786 1297 2010 1357
rect 2044 1297 2268 1357
rect 2302 1297 2308 1357
rect 1488 1285 2308 1297
rect 2500 1295 2515 1370
rect 2570 1295 2590 1370
rect 2500 1285 2590 1295
rect 2730 1357 2870 1370
rect 2730 1297 2784 1357
rect 2818 1297 2870 1357
rect 894 1250 1380 1260
rect 894 1130 950 1250
rect 1370 1130 1380 1250
rect 894 1120 1380 1130
rect 1490 1200 2304 1285
rect 2730 1200 2870 1297
rect 3015 1357 3105 1390
rect 3860 1370 4630 1407
rect 3015 1297 3042 1357
rect 3076 1297 3105 1357
rect 3015 1280 3105 1297
rect 3250 1357 3390 1370
rect 3250 1297 3300 1357
rect 3334 1297 3390 1357
rect 3250 1200 3390 1297
rect 3535 1295 3545 1370
rect 3600 1295 3610 1370
rect 3535 1285 3610 1295
rect 3810 1357 4630 1370
rect 3810 1297 3816 1357
rect 3850 1297 4074 1357
rect 4108 1297 4332 1357
rect 4366 1297 4590 1357
rect 4624 1297 4630 1357
rect 3810 1200 4630 1297
rect 1490 1180 4630 1200
rect 1490 1110 1510 1180
rect 4610 1110 4630 1180
rect 1490 1090 4630 1110
rect 4820 820 4930 2620
rect 20 800 4930 820
rect 20 750 1450 800
rect 4660 750 4930 800
rect 4970 710 5020 2730
rect -80 640 1450 710
rect 4660 640 5020 710
rect -80 620 5020 640
rect 5120 520 5200 2920
rect -240 420 5200 520
rect 5240 380 5320 3060
rect 6840 3060 7460 3140
rect 6840 2960 6940 3060
rect 7360 2960 7460 3060
rect 7840 2960 8680 3000
rect 6700 2940 6960 2960
rect 5580 2780 5840 2800
rect 5580 2300 5600 2780
rect 5820 2300 5840 2780
rect 6700 2760 6720 2940
rect 6940 2760 6960 2940
rect 7340 2940 7600 2960
rect 6700 2749 6877 2760
rect 6911 2749 6960 2760
rect 6700 2740 6960 2749
rect 7129 2925 7175 2937
rect 7129 2749 7135 2925
rect 7169 2749 7175 2925
rect 6871 2737 6917 2740
rect 7129 2737 7175 2749
rect 7340 2760 7360 2940
rect 7580 2760 7600 2940
rect 7340 2749 7393 2760
rect 7427 2749 7600 2760
rect 7340 2740 7600 2749
rect 7640 2940 8380 2960
rect 7640 2760 7660 2940
rect 7760 2760 8380 2940
rect 7640 2740 8380 2760
rect 8460 2740 8680 2960
rect 7387 2737 7433 2740
rect 6927 2700 7119 2705
rect 7185 2700 7377 2705
rect 7840 2700 8680 2740
rect 6920 2699 7380 2700
rect 6920 2665 6939 2699
rect 7107 2665 7197 2699
rect 7365 2665 7380 2699
rect 6920 2600 7380 2665
rect 6920 2420 6940 2600
rect 7360 2420 7380 2600
rect 6920 2400 7380 2420
rect 5580 2280 5840 2300
rect 6920 2300 7380 2320
rect 6920 2120 6940 2300
rect 7360 2120 7380 2300
rect 6920 2054 7380 2120
rect 6920 2020 6939 2054
rect 7107 2020 7197 2054
rect 7365 2020 7380 2054
rect 6927 2014 7119 2020
rect 7185 2014 7377 2020
rect 7840 1980 8680 2020
rect 6700 1961 6960 1980
rect 6700 1960 6877 1961
rect 6911 1960 6960 1961
rect 6700 1780 6720 1960
rect 6940 1780 6960 1960
rect 6700 1760 6960 1780
rect 7100 1961 7200 1980
rect 7100 1785 7135 1961
rect 7169 1785 7200 1961
rect 7100 1680 7200 1785
rect 7340 1961 7600 1980
rect 7340 1960 7393 1961
rect 7427 1960 7600 1961
rect 7340 1780 7360 1960
rect 7580 1780 7600 1960
rect 7340 1760 7600 1780
rect 7640 1960 8680 1980
rect 7640 1780 7660 1960
rect 7760 1780 8560 1960
rect 7640 1760 8560 1780
rect 7840 1740 8560 1760
rect 8640 1740 8680 1960
rect 7840 1720 8680 1740
rect 6840 1600 7460 1680
rect 6840 1500 6940 1600
rect 7360 1500 7460 1600
rect 7840 1500 8680 1540
rect 6700 1480 6960 1500
rect 6700 1300 6720 1480
rect 6940 1300 6960 1480
rect 7340 1480 7600 1500
rect 6700 1289 6877 1300
rect 6911 1289 6960 1300
rect 6700 1280 6960 1289
rect 7129 1465 7175 1477
rect 7129 1289 7135 1465
rect 7169 1289 7175 1465
rect 6871 1277 6917 1280
rect 7129 1277 7175 1289
rect 7340 1300 7360 1480
rect 7580 1300 7600 1480
rect 7340 1289 7393 1300
rect 7427 1289 7600 1300
rect 7340 1280 7600 1289
rect 7640 1480 8380 1500
rect 7640 1300 7660 1480
rect 7760 1300 8380 1480
rect 7640 1280 8380 1300
rect 8460 1280 8680 1500
rect 7387 1277 7433 1280
rect 6927 1240 7119 1245
rect 7185 1240 7377 1245
rect 7840 1240 8680 1280
rect 6920 1239 7380 1240
rect 6920 1205 6939 1239
rect 7107 1205 7197 1239
rect 7365 1205 7380 1239
rect 5420 1180 5560 1200
rect 5420 740 5440 1180
rect 5540 740 5560 1180
rect 6920 1140 7380 1205
rect 6920 960 6940 1140
rect 7360 960 7380 1140
rect 6920 940 7380 960
rect 5420 720 5560 740
rect 6558 600 7570 620
rect 6558 540 6580 600
rect 7540 589 7570 600
rect 7541 555 7570 589
rect 7540 540 7570 555
rect 6558 524 7570 540
rect -380 320 5320 380
rect 6200 360 7200 380
rect 5600 321 5800 340
rect 5600 320 5682 321
rect 5720 320 5800 321
rect 3520 198 4680 200
rect 3516 180 4680 198
rect 3516 100 3540 180
rect 4660 100 4680 180
rect 3516 80 4680 100
rect 3516 -40 4104 80
rect 5600 60 5620 320
rect 3516 -78 3644 -40
rect 4041 -78 4104 -40
rect 3516 -114 4104 -78
rect 4820 40 5620 60
rect 4820 -140 4840 40
rect 5780 -140 5800 320
rect 6200 180 6220 360
rect 6400 284 7200 360
rect 6400 250 6702 284
rect 7190 250 7200 284
rect 6400 180 7200 250
rect 6200 160 7200 180
rect 7300 360 7700 380
rect 7300 348 7500 360
rect 7300 184 7314 348
rect 7362 184 7500 348
rect 7300 180 7500 184
rect 7680 180 7700 360
rect 7300 160 7700 180
rect 6558 60 7570 76
rect 6558 0 6580 60
rect 7560 0 7570 60
rect 6558 -20 7570 0
rect 4820 -160 5800 -140
<< via1 >>
rect 6940 3580 7360 3760
rect 6720 3245 6877 3420
rect 6877 3245 6911 3420
rect 6911 3245 6940 3420
rect 6720 3240 6940 3245
rect 7360 3245 7393 3420
rect 7393 3245 7427 3420
rect 7427 3245 7580 3420
rect 7360 3240 7580 3245
rect 8560 3200 8640 3420
rect 1450 3060 4660 3100
rect 1450 3020 4660 3060
rect 1450 2940 4660 3020
rect 1450 2360 4610 2380
rect 1450 2320 4580 2360
rect 4580 2320 4610 2360
rect 1450 2300 4610 2320
rect 1710 2050 1752 2110
rect 1752 2050 1786 2110
rect 1786 2050 1820 2110
rect 2230 2050 2268 2110
rect 2268 2050 2302 2110
rect 2302 2050 2340 2110
rect 2740 2044 2784 2110
rect 2784 2044 2818 2110
rect 2818 2044 2850 2110
rect 2740 2000 2850 2044
rect 3260 2050 3300 2120
rect 3300 2050 3334 2120
rect 3334 2050 3370 2120
rect 3780 2044 3816 2120
rect 3816 2044 3850 2120
rect 3850 2044 3890 2120
rect 3780 2000 3890 2044
rect 4290 2050 4332 2120
rect 4332 2050 4366 2120
rect 4366 2050 4400 2120
rect 1710 1730 1752 1790
rect 1752 1730 1786 1790
rect 1786 1730 1820 1790
rect 2090 1740 2180 1900
rect 2230 1730 2268 1790
rect 2268 1730 2302 1790
rect 2302 1730 2340 1790
rect 1970 1620 2010 1680
rect 2010 1620 2044 1680
rect 2044 1620 2080 1680
rect 2490 1620 2526 1680
rect 2526 1620 2560 1680
rect 2560 1620 2600 1680
rect 2740 1730 2784 1790
rect 2784 1730 2818 1790
rect 2818 1730 2850 1790
rect 3010 1620 3042 1680
rect 3042 1620 3076 1680
rect 3076 1620 3120 1680
rect 3260 1730 3300 1790
rect 3300 1730 3334 1790
rect 3334 1730 3370 1790
rect 3520 1620 3558 1680
rect 3558 1620 3592 1680
rect 3592 1620 3630 1680
rect 3780 1730 3816 1790
rect 3816 1730 3850 1790
rect 3850 1730 3890 1790
rect 4160 1750 4240 1900
rect 4030 1620 4074 1680
rect 4074 1620 4108 1680
rect 4108 1620 4140 1680
rect 4290 1730 4332 1790
rect 4332 1730 4366 1790
rect 4366 1730 4400 1790
rect 2950 1441 3170 1490
rect 2950 1430 3014 1441
rect 3014 1430 3104 1441
rect 3104 1430 3170 1441
rect 2515 1357 2570 1370
rect 2515 1297 2526 1357
rect 2526 1297 2560 1357
rect 2560 1297 2570 1357
rect 2515 1295 2570 1297
rect 950 1230 1370 1250
rect 950 1140 960 1230
rect 960 1140 1360 1230
rect 1360 1140 1370 1230
rect 950 1130 1370 1140
rect 3545 1357 3600 1370
rect 3545 1297 3558 1357
rect 3558 1297 3592 1357
rect 3592 1297 3600 1357
rect 3545 1295 3600 1297
rect 1510 1170 4610 1180
rect 1510 1120 1530 1170
rect 1530 1120 4580 1170
rect 4580 1120 4610 1170
rect 1510 1110 4610 1120
rect 1450 750 4660 800
rect 1450 710 4660 750
rect 1450 640 4660 710
rect 5600 2720 5820 2780
rect 5600 2320 5640 2720
rect 5640 2320 5760 2720
rect 5760 2320 5820 2720
rect 5600 2300 5820 2320
rect 6720 2925 6940 2940
rect 6720 2760 6877 2925
rect 6877 2760 6911 2925
rect 6911 2760 6940 2925
rect 7360 2925 7580 2940
rect 7360 2760 7393 2925
rect 7393 2760 7427 2925
rect 7427 2760 7580 2925
rect 8380 2740 8460 2960
rect 6940 2420 7360 2600
rect 6940 2120 7360 2300
rect 6720 1785 6877 1960
rect 6877 1785 6911 1960
rect 6911 1785 6940 1960
rect 6720 1780 6940 1785
rect 7360 1785 7393 1960
rect 7393 1785 7427 1960
rect 7427 1785 7580 1960
rect 7360 1780 7580 1785
rect 8560 1740 8640 1960
rect 6720 1465 6940 1480
rect 6720 1300 6877 1465
rect 6877 1300 6911 1465
rect 6911 1300 6940 1465
rect 7360 1465 7580 1480
rect 7360 1300 7393 1465
rect 7393 1300 7427 1465
rect 7427 1300 7580 1465
rect 8380 1280 8460 1500
rect 5440 740 5540 1180
rect 6940 960 7360 1140
rect 6580 589 7540 600
rect 6580 555 6587 589
rect 6587 555 6621 589
rect 6621 555 6679 589
rect 6679 555 6713 589
rect 6713 555 6771 589
rect 6771 555 6805 589
rect 6805 555 6863 589
rect 6863 555 6897 589
rect 6897 555 6955 589
rect 6955 555 6989 589
rect 6989 555 7047 589
rect 7047 555 7081 589
rect 7081 555 7139 589
rect 7139 555 7173 589
rect 7173 555 7231 589
rect 7231 555 7265 589
rect 7265 555 7323 589
rect 7323 555 7357 589
rect 7357 555 7415 589
rect 7415 555 7449 589
rect 7449 555 7507 589
rect 7507 555 7540 589
rect 6580 540 7540 555
rect 3540 100 4660 180
rect 5620 40 5682 320
rect 4840 -40 5682 40
rect 4840 -78 4843 -40
rect 4843 -78 5240 -40
rect 5240 -76 5682 -40
rect 5682 -76 5720 320
rect 5720 -76 5780 320
rect 5240 -78 5780 -76
rect 4840 -140 5780 -78
rect 6220 180 6400 360
rect 7500 180 7680 360
rect 6580 45 7560 60
rect 6580 11 6587 45
rect 6587 11 6621 45
rect 6621 11 6679 45
rect 6679 11 6713 45
rect 6713 11 6771 45
rect 6771 11 6805 45
rect 6805 11 6863 45
rect 6863 11 6897 45
rect 6897 11 6955 45
rect 6955 11 6989 45
rect 6989 11 7047 45
rect 7047 11 7081 45
rect 7081 11 7139 45
rect 7139 11 7173 45
rect 7173 11 7231 45
rect 7231 11 7265 45
rect 7265 11 7323 45
rect 7323 11 7357 45
rect 7357 11 7415 45
rect 7415 11 7449 45
rect 7449 11 7507 45
rect 7507 11 7541 45
rect 7541 11 7560 45
rect 6580 0 7560 11
<< metal2 >>
rect 6400 3760 7780 3780
rect 6400 3580 6540 3760
rect 6860 3580 6940 3760
rect 7360 3580 7780 3760
rect 6400 3560 7780 3580
rect -840 3420 7780 3440
rect -840 3240 -820 3420
rect -520 3240 6720 3420
rect 6940 3240 7360 3420
rect 7580 3240 7780 3420
rect -840 3220 7780 3240
rect 8540 3420 8660 3440
rect 8540 3200 8560 3420
rect 8640 3200 8660 3420
rect 8540 3180 8660 3200
rect 1430 3100 4680 3120
rect 1430 2940 1450 3100
rect 4660 2940 4680 3100
rect 8360 2960 8480 2980
rect 1430 2540 4680 2940
rect 6400 2940 8280 2960
rect 1430 2270 1440 2540
rect 4670 2270 4680 2540
rect 5580 2780 5840 2800
rect 5580 2300 5600 2780
rect 5820 2300 5840 2780
rect 6400 2760 6720 2940
rect 6940 2760 7360 2940
rect 7580 2760 7980 2940
rect 8260 2760 8280 2940
rect 6400 2740 8280 2760
rect 8360 2740 8380 2960
rect 8460 2740 8480 2960
rect 8360 2720 8480 2740
rect 5580 2280 5840 2300
rect 6400 2600 7780 2620
rect 6400 2420 6940 2600
rect 7360 2420 7500 2600
rect 6400 2300 7500 2420
rect 1430 2260 4680 2270
rect 1700 2110 1830 2120
rect 1700 2050 1710 2110
rect 1820 2050 1830 2110
rect 1700 1800 1830 2050
rect 1700 1730 1710 1800
rect 1820 1730 1830 1800
rect 1700 1720 1830 1730
rect 1860 2110 2190 2120
rect 1860 1890 1870 2110
rect 2140 1900 2190 2110
rect 1860 1740 2090 1890
rect 2180 1740 2190 1900
rect 1860 1720 2190 1740
rect 2220 2110 2350 2120
rect 2220 2040 2230 2110
rect 2340 2040 2350 2110
rect 2220 1790 2350 2040
rect 2220 1730 2230 1790
rect 2340 1730 2350 1790
rect 2220 1720 2350 1730
rect 2730 2110 2860 2130
rect 2730 2000 2740 2110
rect 2850 2000 2860 2110
rect 2730 1800 2860 2000
rect 2730 1730 2740 1800
rect 2850 1730 2860 1800
rect 2730 1720 2860 1730
rect 3250 2120 3380 2130
rect 3250 2040 3260 2120
rect 3370 2040 3380 2120
rect 3250 1790 3380 2040
rect 3250 1730 3260 1790
rect 3370 1730 3380 1790
rect 3250 1720 3380 1730
rect 3770 2120 3900 2130
rect 3770 2000 3780 2120
rect 3890 2000 3900 2120
rect 3770 1800 3900 2000
rect 4280 2120 4410 2130
rect 4280 2040 4290 2120
rect 4400 2040 4410 2120
rect 6400 2120 6940 2300
rect 7360 2120 7500 2300
rect 7680 2120 7780 2600
rect 6400 2100 7780 2120
rect 3770 1730 3780 1800
rect 3890 1730 3900 1800
rect 3950 1910 4250 1920
rect 3950 1740 3970 1910
rect 4240 1740 4250 1910
rect 3950 1730 4250 1740
rect 4280 1790 4410 2040
rect 4280 1730 4290 1790
rect 4400 1730 4410 1790
rect 5940 1960 7780 1980
rect 5940 1780 5960 1960
rect 6160 1780 6720 1960
rect 6940 1780 7360 1960
rect 7580 1780 7780 1960
rect 5940 1760 7780 1780
rect 8540 1960 8660 1980
rect 3770 1720 3900 1730
rect 4280 1720 4410 1730
rect 8540 1740 8560 1960
rect 8640 1740 8660 1960
rect 8540 1720 8660 1740
rect 1950 1680 4160 1690
rect 1950 1620 1970 1680
rect 2080 1620 2490 1680
rect 2600 1620 3010 1680
rect 3120 1620 3520 1680
rect 3630 1620 4030 1680
rect 4140 1620 4160 1680
rect 1950 1600 4160 1620
rect 940 1490 3200 1530
rect 940 1430 2950 1490
rect 3170 1430 3200 1490
rect 940 1420 3200 1430
rect 940 1250 1380 1420
rect 3270 1385 3630 1600
rect 8360 1500 8480 1520
rect 2480 1370 3630 1385
rect 2480 1295 2515 1370
rect 2570 1295 3545 1370
rect 3600 1295 3630 1370
rect 2480 1280 3630 1295
rect 6400 1480 8280 1500
rect 6400 1300 6720 1480
rect 6940 1300 7360 1480
rect 7580 1300 7980 1480
rect 8260 1300 8280 1480
rect 6400 1280 8280 1300
rect 8360 1280 8380 1500
rect 8460 1280 8480 1500
rect 8360 1260 8480 1280
rect 940 1130 950 1250
rect 1370 1130 1380 1250
rect 940 1120 1380 1130
rect 1430 970 1450 1220
rect 4660 1180 5580 1220
rect 4660 970 5440 1180
rect 1430 800 5440 970
rect 1430 640 1450 800
rect 4660 740 5440 800
rect 5540 740 5580 1180
rect 6400 1140 7780 1160
rect 6400 960 6460 1140
rect 6860 960 6940 1140
rect 7360 960 7780 1140
rect 6400 940 7780 960
rect 4660 700 5580 740
rect 6460 700 7580 720
rect 4660 640 4680 700
rect 1430 620 4680 640
rect 3520 180 4680 620
rect 6460 600 6980 700
rect 7360 600 7580 700
rect 6460 540 6580 600
rect 7540 540 7580 600
rect 6460 520 7580 540
rect 6200 360 6420 380
rect 3520 100 3540 180
rect 4660 100 4680 180
rect 3520 60 4680 100
rect 5600 320 5800 340
rect 5600 60 5620 320
rect 4820 40 5620 60
rect 4820 -140 4840 40
rect 5780 -140 5800 320
rect 6200 180 6220 360
rect 6400 180 6420 360
rect 6200 160 6420 180
rect 7480 360 7700 380
rect 7480 180 7500 360
rect 7680 180 7700 360
rect 7480 160 7700 180
rect 6460 60 7580 80
rect 6460 -100 6540 60
rect 7560 0 7580 60
rect 6860 -100 7580 0
rect 6460 -120 7580 -100
rect 4820 -160 5800 -140
<< via2 >>
rect 6540 3580 6860 3760
rect -820 3240 -520 3420
rect 8560 3200 8640 3420
rect 1440 2380 4670 2540
rect 1440 2300 1450 2380
rect 1450 2300 4610 2380
rect 4610 2300 4670 2380
rect 1440 2270 4670 2300
rect 5600 2300 5820 2780
rect 7980 2760 8260 2940
rect 8380 2740 8460 2960
rect 1710 1790 1820 1800
rect 1710 1730 1820 1790
rect 1870 1900 2140 2110
rect 1870 1890 2090 1900
rect 2090 1890 2140 1900
rect 2230 2050 2340 2110
rect 2230 2040 2340 2050
rect 2740 1790 2850 1800
rect 2740 1730 2850 1790
rect 3260 2050 3370 2110
rect 3260 2040 3370 2050
rect 4290 2050 4400 2110
rect 4290 2040 4400 2050
rect 7500 2120 7680 2600
rect 3780 1790 3890 1800
rect 3780 1730 3890 1790
rect 3970 1900 4240 1910
rect 3970 1750 4160 1900
rect 4160 1750 4240 1900
rect 3970 1740 4240 1750
rect 5960 1780 6160 1960
rect 8560 1740 8640 1960
rect 7980 1300 8260 1480
rect 8380 1280 8460 1500
rect 1450 1180 4660 1220
rect 1450 1110 1510 1180
rect 1510 1110 4610 1180
rect 4610 1110 4660 1180
rect 1450 970 4660 1110
rect 6460 960 6860 1140
rect 6980 600 7360 700
rect 6980 540 7360 600
rect 5620 40 5780 320
rect 4840 -140 5780 40
rect 6220 180 6400 360
rect 7500 180 7680 360
rect 6540 0 6580 60
rect 6580 0 6860 60
rect 6540 -100 6860 0
<< metal3 >>
rect -840 3420 -500 4140
rect -840 3240 -820 3420
rect -520 3240 -500 3420
rect -840 2180 -500 3240
rect 6520 3760 6880 4280
rect 6520 3580 6540 3760
rect 6860 3580 6880 3760
rect -380 3060 5320 3120
rect -380 2320 -320 3060
rect 5240 2320 5320 3060
rect -380 2270 1440 2320
rect 4670 2270 5320 2320
rect -380 2260 5320 2270
rect 5580 2780 5840 2800
rect 5580 2300 5600 2780
rect 5820 2300 5840 2780
rect 5580 2240 5840 2300
rect -840 2110 2150 2180
rect 5580 2140 6180 2240
rect 4040 2120 6180 2140
rect -840 1890 1870 2110
rect 2140 1890 2150 2110
rect -840 1880 2150 1890
rect 1480 1870 2150 1880
rect 2210 2110 6180 2120
rect 2210 2040 2230 2110
rect 2340 2040 3260 2110
rect 3370 2040 4290 2110
rect 4400 2040 6180 2110
rect 2210 2030 4410 2040
rect 2210 1870 3870 2030
rect 3960 1960 4630 1970
rect 5940 1960 6180 2040
rect 3960 1910 5800 1960
rect 1700 1800 3900 1810
rect 1700 1730 1710 1800
rect 1820 1730 2740 1800
rect 2850 1730 3780 1800
rect 3890 1730 3900 1800
rect 1700 1720 3900 1730
rect 2240 1560 3900 1720
rect 3960 1740 3970 1910
rect 4240 1740 5800 1910
rect 5940 1780 5960 1960
rect 6160 1780 6180 1960
rect 5940 1760 6180 1780
rect 3960 1580 5800 1740
rect -380 1220 5320 1250
rect -380 1200 1450 1220
rect 4660 1200 5320 1220
rect -380 380 -320 1200
rect 5260 380 5320 1200
rect -380 320 5320 380
rect 5600 320 5800 1580
rect 6520 1200 6880 3580
rect 5600 60 5620 320
rect 4820 40 5620 60
rect 4820 -140 4840 40
rect 5780 -140 5800 320
rect 6200 1140 6880 1200
rect 6200 960 6460 1140
rect 6860 960 6880 1140
rect 6200 880 6880 960
rect 6960 3100 7380 3120
rect 6960 2280 6980 3100
rect 7360 2280 7380 3100
rect 7960 2940 8280 4280
rect 8540 3420 8660 3440
rect 8540 3200 8560 3420
rect 8640 3200 8660 3420
rect 8540 3100 8660 3200
rect 7960 2760 7980 2940
rect 8260 2760 8280 2940
rect 6200 360 6420 880
rect 6200 180 6220 360
rect 6400 180 6420 360
rect 6200 160 6420 180
rect 6520 700 6880 720
rect 6520 340 6540 700
rect 6860 340 6880 700
rect 6960 700 7380 2280
rect 6960 540 6980 700
rect 7360 540 7380 700
rect 6960 520 7380 540
rect 7480 2600 7700 2620
rect 7480 2120 7500 2600
rect 7680 2120 7700 2600
rect 6520 60 6880 340
rect 7480 360 7700 2120
rect 7960 1480 8280 2760
rect 7960 1300 7980 1480
rect 8260 1300 8280 1480
rect 7960 1280 8280 1300
rect 8360 2960 8480 2980
rect 8360 2740 8380 2960
rect 8460 2740 8480 2960
rect 8360 1500 8480 2740
rect 8540 2280 8560 3100
rect 8640 2280 8660 3100
rect 8540 1960 8660 2280
rect 8540 1740 8560 1960
rect 8640 1740 8660 1960
rect 8540 1720 8660 1740
rect 8360 1280 8380 1500
rect 8460 1280 8480 1500
rect 7480 180 7500 360
rect 7680 180 7700 360
rect 8360 1240 8480 1280
rect 8360 340 8380 1240
rect 8460 340 8480 1240
rect 8360 320 8480 340
rect 7480 160 7700 180
rect 6520 -100 6540 60
rect 6860 -100 6880 60
rect 6520 -120 6880 -100
rect 4820 -160 5800 -140
<< via3 >>
rect -320 2540 5240 3060
rect -320 2320 1440 2540
rect 1440 2320 4670 2540
rect 4670 2320 5240 2540
rect -320 970 1450 1200
rect 1450 970 4660 1200
rect 4660 970 5260 1200
rect -320 380 5260 970
rect 6980 2280 7360 3100
rect 6540 340 6860 700
rect 8560 2280 8640 3100
rect 8380 340 8460 1240
<< metal4 >>
rect -380 3100 9200 3120
rect -380 3060 6980 3100
rect -380 2320 -320 3060
rect 5240 2320 6980 3060
rect -380 2280 6980 2320
rect 7360 2280 8560 3100
rect 8640 2280 9200 3100
rect -380 2260 9200 2280
rect -380 1240 9200 1260
rect -380 1200 8380 1240
rect -380 380 -320 1200
rect 5260 700 8380 1200
rect 5260 380 6540 700
rect -380 340 6540 380
rect 6860 340 8380 700
rect 8460 340 9200 1240
rect -380 320 9200 340
<< labels >>
flabel metal3 6520 3760 6880 4280 0 FreeSans 1600 0 0 0 CTRL
port 2 nsew
flabel via3 -320 380 5260 1200 0 FreeSans 1600 0 0 0 VSS
port 5 nsew
flabel via3 -320 2320 5240 3060 0 FreeSans 1600 0 0 0 VDD
port 4 nsew
flabel metal3 7960 2940 8280 4280 0 FreeSans 1600 0 0 0 OUT
port 3 nsew
flabel metal3 -840 3420 -500 4140 0 FreeSans 1600 0 0 0 IN
port 1 nsew
flabel metal2 6400 1760 6720 1980 0 FreeSans 1600 0 0 0 tgate_1.IN
flabel metal2 6400 1280 6720 1500 0 FreeSans 1600 0 0 0 tgate_1.OUT
flabel metal2 6400 2100 6940 2320 0 FreeSans 1600 0 0 0 tgate_1.CTRLB
flabel metal2 6400 940 6940 1160 0 FreeSans 1600 0 0 0 tgate_1.CTRL
flabel metal1 7760 1760 8080 1980 0 FreeSans 1600 0 0 0 tgate_1.VDD
flabel metal1 7760 1280 8080 1500 0 FreeSans 1600 0 0 0 tgate_1.VSS
flabel metal2 6400 3220 6720 3440 0 FreeSans 1600 0 0 0 tgate_0.IN
flabel metal2 6400 2740 6720 2960 0 FreeSans 1600 0 0 0 tgate_0.OUT
flabel metal2 6400 3560 6940 3780 0 FreeSans 1600 0 0 0 tgate_0.CTRLB
flabel metal2 6400 2400 6940 2620 0 FreeSans 1600 0 0 0 tgate_0.CTRL
flabel metal1 7760 3220 8080 3440 0 FreeSans 1600 0 0 0 tgate_0.VDD
flabel metal1 7760 2740 8080 2960 0 FreeSans 1600 0 0 0 tgate_0.VSS
flabel metal1 7405 14 7453 40 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tap_2_0.VGND
flabel metal1 7407 561 7461 583 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tap_2_0.VPWR
flabel locali 7421 459 7446 484 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__tap_2_0.VPB
flabel locali 7506 120 7541 150 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__tap_2_0.VNB
flabel locali 7514 453 7536 482 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__tap_2_0.VPB
rlabel comment 7386 28 7386 28 4 sky130_fd_sc_hd__tap_2_0.tap_2
rlabel metal1 7386 -20 7570 76 1 sky130_fd_sc_hd__tap_2_0.VGND
rlabel metal1 7386 524 7570 620 1 sky130_fd_sc_hd__tap_2_0.VPWR
flabel locali 6771 249 6805 283 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__inv_8_0.A
flabel locali 6863 249 6897 283 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__inv_8_0.A
flabel locali 6955 249 6989 283 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__inv_8_0.A
flabel locali 7047 249 7081 283 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__inv_8_0.A
flabel locali 7139 249 7173 283 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__inv_8_0.A
flabel locali 7231 249 7265 283 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__inv_8_0.A
flabel locali 7323 249 7357 283 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__inv_8_0.Y
flabel locali 6587 249 6621 283 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__inv_8_0.Y
flabel pwell 6587 11 6621 45 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_8_0.VNB
flabel nwell 6587 555 6621 589 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_8_0.VPB
flabel metal1 6587 11 6621 45 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_8_0.VGND
flabel metal1 6587 555 6621 589 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_8_0.VPWR
rlabel comment 6558 28 6558 28 4 sky130_fd_sc_hd__inv_8_0.inv_8
rlabel metal1 6558 -20 7386 76 1 sky130_fd_sc_hd__inv_8_0.VGND
rlabel metal1 6558 524 7386 620 1 sky130_fd_sc_hd__inv_8_0.VPWR
flabel metal3 4240 1580 4630 1970 0 FreeSans 800 0 0 0 myOpamp_0.INn
flabel metal3 2210 1870 3870 2120 0 FreeSans 800 0 0 0 myOpamp_0.OUT
flabel metal3 1450 970 4660 1220 0 FreeSans 800 0 0 0 myOpamp_0.VSS
flabel metal3 1440 2270 4670 2540 0 FreeSans 800 0 0 0 myOpamp_0.VDD
flabel metal3 1480 1870 1870 2180 0 FreeSans 800 0 0 0 myOpamp_0.INp
<< end >>
