magic
tech sky130A
magscale 1 2
timestamp 1713227210
<< nmos >>
rect -745 -81 -545 19
rect -487 -81 -287 19
rect -229 -81 -29 19
rect 29 -81 229 19
rect 287 -81 487 19
rect 545 -81 745 19
<< ndiff >>
rect -803 7 -745 19
rect -803 -69 -791 7
rect -757 -69 -745 7
rect -803 -81 -745 -69
rect -545 7 -487 19
rect -545 -69 -533 7
rect -499 -69 -487 7
rect -545 -81 -487 -69
rect -287 7 -229 19
rect -287 -69 -275 7
rect -241 -69 -229 7
rect -287 -81 -229 -69
rect -29 7 29 19
rect -29 -69 -17 7
rect 17 -69 29 7
rect -29 -81 29 -69
rect 229 7 287 19
rect 229 -69 241 7
rect 275 -69 287 7
rect 229 -81 287 -69
rect 487 7 545 19
rect 487 -69 499 7
rect 533 -69 545 7
rect 487 -81 545 -69
rect 745 7 803 19
rect 745 -69 757 7
rect 791 -69 803 7
rect 745 -81 803 -69
<< ndiffc >>
rect -791 -69 -757 7
rect -533 -69 -499 7
rect -275 -69 -241 7
rect -17 -69 17 7
rect 241 -69 275 7
rect 499 -69 533 7
rect 757 -69 791 7
<< poly >>
rect -745 91 -545 107
rect -745 57 -729 91
rect -561 57 -545 91
rect -745 19 -545 57
rect -487 91 -287 107
rect -487 57 -471 91
rect -303 57 -287 91
rect -487 19 -287 57
rect -229 91 -29 107
rect -229 57 -213 91
rect -45 57 -29 91
rect -229 19 -29 57
rect 29 91 229 107
rect 29 57 45 91
rect 213 57 229 91
rect 29 19 229 57
rect 287 91 487 107
rect 287 57 303 91
rect 471 57 487 91
rect 287 19 487 57
rect 545 91 745 107
rect 545 57 561 91
rect 729 57 745 91
rect 545 19 745 57
rect -745 -107 -545 -81
rect -487 -107 -287 -81
rect -229 -107 -29 -81
rect 29 -107 229 -81
rect 287 -107 487 -81
rect 545 -107 745 -81
<< polycont >>
rect -729 57 -561 91
rect -471 57 -303 91
rect -213 57 -45 91
rect 45 57 213 91
rect 303 57 471 91
rect 561 57 729 91
<< locali >>
rect -745 57 -729 91
rect -561 57 -545 91
rect -487 57 -471 91
rect -303 57 -287 91
rect -229 57 -213 91
rect -45 57 -29 91
rect 29 57 45 91
rect 213 57 229 91
rect 287 57 303 91
rect 471 57 487 91
rect 545 57 561 91
rect 729 57 745 91
rect -791 7 -757 23
rect -791 -85 -757 -69
rect -533 7 -499 23
rect -533 -85 -499 -69
rect -275 7 -241 23
rect -275 -85 -241 -69
rect -17 7 17 23
rect -17 -85 17 -69
rect 241 7 275 23
rect 241 -85 275 -69
rect 499 7 533 23
rect 499 -85 533 -69
rect 757 7 791 23
rect 757 -85 791 -69
<< viali >>
rect -729 57 -561 91
rect -471 57 -303 91
rect -213 57 -45 91
rect 45 57 213 91
rect 303 57 471 91
rect 561 57 729 91
rect -791 -69 -757 7
rect -533 -69 -499 7
rect -275 -69 -241 7
rect -17 -69 17 7
rect 241 -69 275 7
rect 499 -69 533 7
rect 757 -69 791 7
<< metal1 >>
rect -741 91 -549 97
rect -741 57 -729 91
rect -561 57 -549 91
rect -741 51 -549 57
rect -483 91 -291 97
rect -483 57 -471 91
rect -303 57 -291 91
rect -483 51 -291 57
rect -225 91 -33 97
rect -225 57 -213 91
rect -45 57 -33 91
rect -225 51 -33 57
rect 33 91 225 97
rect 33 57 45 91
rect 213 57 225 91
rect 33 51 225 57
rect 291 91 483 97
rect 291 57 303 91
rect 471 57 483 91
rect 291 51 483 57
rect 549 91 741 97
rect 549 57 561 91
rect 729 57 741 91
rect 549 51 741 57
rect -797 7 -751 19
rect -797 -69 -791 7
rect -757 -69 -751 7
rect -797 -81 -751 -69
rect -539 7 -493 19
rect -539 -69 -533 7
rect -499 -69 -493 7
rect -539 -81 -493 -69
rect -281 7 -235 19
rect -281 -69 -275 7
rect -241 -69 -235 7
rect -281 -81 -235 -69
rect -23 7 23 19
rect -23 -69 -17 7
rect 17 -69 23 7
rect -23 -81 23 -69
rect 235 7 281 19
rect 235 -69 241 7
rect 275 -69 281 7
rect 235 -81 281 -69
rect 493 7 539 19
rect 493 -69 499 7
rect 533 -69 539 7
rect 493 -81 539 -69
rect 751 7 797 19
rect 751 -69 757 7
rect 791 -69 797 7
rect 751 -81 797 -69
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.5 l 1 m 1 nf 6 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
