* NGSPICE file created from guitpedal_flat.ext - technology: sky130A

.subckt tt_um_guitar_pedal ua[0] ua[1] ui_in[0] VPWR ui_in[1] VGND ui_in[2] ui_in[3] ui_in[4] ui_in[5]
+ ui_in[6] ui_in[7]
X0 VGND.t245 ui_in[4].t0 distortionUnit_5.tgate_1.CTRLB VGND.t244 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_20524_36601# a_20524_36601# VPWR.t212 VPWR.t211 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2 VGND.t406 VGND.t405 VGND.t406 VGND.t134 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X3 distortionUnit_0.tgate_1.CTRLB ui_in[6].t0 VPWR.t271 distortionUnit_0.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR.t270 VPWR.t268 distortionUnit_0.tgate_1.IN VPWR.t269 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X5 a_7876_23853# VGND.t403 VGND.t404 VGND.t331 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X6 VGND.t402 VGND.t400 VGND.t402 VGND.t401 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X7 VPWR.t49 a_7752_16807# a_7752_16807# VPWR.t48 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X8 distortionUnit_4.IN ui_in[3].t0 distortionUnit_5.IN.t3 VPWR.t133 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X9 ua[1].t5 ui_in[7].t0 distortionUnit_7.IN VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X10 distortionUnit_6.IN ui_in[4].t1 distortionUnit_5.tgate_1.IN VGND.t243 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X11 ua[0].t3 distortionUnit_1.tgate_1.CTRLB distortionUnit_2.IN VGND.t204 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X12 a_7752_16807# distortionUnit_6.OUT a_8010_16807# VGND.t46 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X13 distortionUnit_4.tgate_1.IN distortionUnit_4.myOpamp_0.INn a_20746_30481# VGND.t100 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X14 VPWR.t129 a_20934_16677# distortionUnit_7.tgate_1.IN VPWR.t128 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X15 ua[1].t1 distortionUnit_7.tgate_1.CTRLB distortionUnit_7.IN VGND.t199 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X16 VGND.t399 VGND.t398 VGND.t399 VGND.t211 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X17 distortionUnit_1.tgate_1.IN distortionUnit_1.myOpamp_0.INn a_7968_36445# VGND.t56 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X18 distortionUnit_7.tgate_1.IN distortionUnit_7.myOpamp_0.INn a_21192_16677# VGND.t324 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X19 a_7752_16807# distortionUnit_6.OUT a_8010_16807# VGND.t44 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X20 VPWR.t89 ui_in[2].t0 distortionUnit_3.tgate_1.CTRLB distortionUnit_3.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 distortionUnit_2.IN distortionUnit_1.tgate_1.CTRLB distortionUnit_1.tgate_1.IN VPWR.t181 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X22 VPWR.t185 ui_in[6].t1 distortionUnit_0.tgate_1.CTRLB distortionUnit_0.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X23 distortionUnit_6.tgate_1.CTRLB ui_in[5].t0 VPWR.t78 distortionUnit_6.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 VGND.t144 a_19680_36146# a_20782_36601# VGND.t143 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X25 distortionUnit_0.tgate_1.IN a_7752_16807# VPWR.t47 VPWR.t46 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X26 VGND.t182 ui_in[3].t1 distortionUnit_4.tgate_1.CTRLB VGND.t181 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X27 distortionUnit_4.tgate_1.CTRLB ui_in[3].t2 VGND.t4 VGND.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X28 a_20782_36601# distortionUnit_2.myOpamp_0.INn distortionUnit_2.tgate_1.IN VGND.t135 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X29 VPWR.t2 ui_in[6].t2 distortionUnit_0.tgate_1.CTRLB distortionUnit_0.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 VGND.t130 a_19644_30026# a_20746_30481# VGND.t129 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X31 distortionUnit_7.IN ui_in[6].t3 distortionUnit_6.OUT VPWR.t4 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X32 distortionUnit_7.IN distortionUnit_7.tgate_1.CTRLB ua[1].t0 VGND.t198 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X33 a_7752_16807# VPWR.t265 VPWR.t267 VPWR.t266 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X34 distortionUnit_6.tgate_1.IN ui_in[5].t1 distortionUnit_6.OUT VGND.t438 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X35 distortionUnit_3.tgate_1.CTRLB ui_in[2].t1 VPWR.t12 distortionUnit_3.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X36 a_7876_23853# a_7876_23853# VPWR.t74 VPWR.t73 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X37 VPWR.t264 VPWR.t262 distortionUnit_7.tgate_1.IN VPWR.t263 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X38 a_8010_16807# distortionUnit_0.myOpamp_0.INn distortionUnit_0.tgate_1.IN VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X39 a_20746_30481# distortionUnit_4.IN a_20488_30481# VGND.t321 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X40 VGND.t88 a_6912_30102# a_8014_30557# VGND.t87 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X41 VPWR.t156 a_7756_30557# a_7756_30557# VPWR.t155 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X42 VGND.t459 a_20090_16222# a_21192_16677# VGND.t59 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X43 distortionUnit_3.tgate_1.CTRLB ui_in[2].t2 VPWR.t1 distortionUnit_3.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X44 VGND.t397 VGND.t396 distortionUnit_3.tgate_1.IN VGND.t316 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X45 distortionUnit_5.tgate_1.CTRLB ui_in[4].t2 VGND.t242 VGND.t241 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X46 distortionUnit_6.tgate_1.IN distortionUnit_6.myOpamp_0.INn a_20842_23723# VGND.t32 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X47 VPWR.t261 VPWR.t259 distortionUnit_2.tgate_1.IN VPWR.t260 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X48 distortionUnit_0.tgate_1.CTRLB ui_in[6].t4 VPWR.t10 distortionUnit_0.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X49 a_9762_22154# distortionUnit_5.myOpamp_0.INn VGND.t424 sky130_fd_pr__res_xhigh_po_0p35 l=4
X50 a_8134_23853# distortionUnit_5.myOpamp_0.INn distortionUnit_5.tgate_1.IN VGND.t163 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X51 a_20782_36601# a_19680_36146# VGND.t142 VGND.t133 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X52 a_8014_30557# distortionUnit_3.IN a_7756_30557# VGND.t81 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X53 VPWR a_19680_36146# VGND sky130_fd_pr__res_xhigh_po_0p35 l=26.11
X54 distortionUnit_4.tgate_1.CTRLB ui_in[3].t3 VGND.t222 VGND.t221 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X55 VGND.t395 VGND.t394 VGND.t395 VGND.t361 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X56 VPWR.t186 a_19740_23268# VGND.t219 sky130_fd_pr__res_xhigh_po_0p35 l=0.16
X57 distortionUnit_5.tgate_1.CTRLB ui_in[4].t3 VGND.t240 VGND.t239 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X58 distortionUnit_6.OUT distortionUnit_0.tgate_1.CTRLB distortionUnit_7.IN VGND.t20 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X59 distortionUnit_2.IN ui_in[1].t0 distortionUnit_3.IN VPWR.t184 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X60 a_6908_16352# a_6908_16352# VGND.t51 VGND.t50 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X61 distortionUnit_1.tgate_1.CTRLB ui_in[0].t0 VPWR.t307 distortionUnit_1.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X62 VPWR.t80 ui_in[0].t1 distortionUnit_1.tgate_1.CTRLB distortionUnit_1.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X63 distortionUnit_7.tgate_1.IN a_20934_16677# VPWR.t127 VPWR.t126 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X64 VGND.t209 ui_in[1].t1 distortionUnit_2.tgate_1.CTRLB VGND.t208 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X65 distortionUnit_4.tgate_1.IN a_20488_30481# VPWR.t179 VPWR.t178 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X66 distortionUnit_6.tgate_1.IN a_20584_23723# VPWR.t296 VPWR.t295 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X67 distortionUnit_2.tgate_1.CTRLB ui_in[1].t2 VGND.t227 VGND.t226 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X68 a_21192_16677# a_20090_16222# VGND.t458 VGND.t434 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X69 a_6866_35990# a_6866_35990# VGND.t451 VGND.t101 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X70 distortionUnit_7.tgate_1.IN a_20934_16677# VPWR.t125 VPWR.t124 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X71 VPWR.t72 a_7876_23853# distortionUnit_5.tgate_1.IN VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X72 distortionUnit_3.tgate_1.IN distortionUnit_3.myOpamp_0.INn a_8014_30557# VGND.t180 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X73 a_20842_23723# distortionUnit_6.IN a_20584_23723# VGND.t214 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X74 a_8014_30557# a_6912_30102# VGND.t86 VGND.t85 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X75 distortionUnit_1.tgate_1.IN ui_in[0].t2 distortionUnit_2.IN VGND.t430 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X76 distortionUnit_5.tgate_1.IN distortionUnit_5.myOpamp_0.INn a_8134_23853# VGND.t159 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X77 a_20842_23723# distortionUnit_6.IN a_20584_23723# VGND.t213 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X78 VGND.t393 VGND.t392 VGND.t393 VGND.t173 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X79 VGND.t391 VGND.t390 VGND.t391 VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X80 VGND.t238 ui_in[4].t4 distortionUnit_5.tgate_1.CTRLB VGND.t237 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X81 distortionUnit_6.tgate_1.CTRLB ui_in[5].t2 VGND.t453 VGND.t452 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X82 distortionUnit_5.tgate_1.IN distortionUnit_5.myOpamp_0.INn a_8134_23853# VGND.t301 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X83 distortionUnit_3.IN ui_in[1].t3 distortionUnit_2.IN VPWR.t25 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X84 VPWR.t54 ui_in[0].t3 distortionUnit_1.tgate_1.CTRLB distortionUnit_1.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X85 a_7756_30557# VGND.t388 VGND.t389 VGND.t297 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X86 distortionUnit_7.tgate_1.IN distortionUnit_7.myOpamp_0.INn VGND.t92 sky130_fd_pr__res_xhigh_po_0p35 l=10
X87 distortionUnit_6.tgate_1.IN distortionUnit_6.tgate_1.CTRLB distortionUnit_6.OUT VPWR.t273 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X88 ua[0].t0 ui_in[0].t4 distortionUnit_2.IN VPWR.t86 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X89 VGND.t387 VGND.t385 VGND.t386 VGND.t352 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0 ps=0 w=0.42 l=1
X90 distortionUnit_4.tgate_1.IN ui_in[3].t4 distortionUnit_5.IN.t1 VGND.t189 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X91 a_20488_30481# distortionUnit_4.IN a_20746_30481# VGND.t123 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X92 VPWR.t123 a_20934_16677# a_20934_16677# VPWR.t122 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X93 distortionUnit_7.tgate_1.CTRLB ui_in[7].t1 VPWR.t24 distortionUnit_7.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X94 VPWR.t177 a_20488_30481# a_20488_30481# VPWR.t176 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X95 VGND.t384 VGND.t383 VGND.t384 VGND.t313 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X96 a_7756_30557# a_7756_30557# VPWR.t154 VPWR.t153 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X97 distortionUnit_2.tgate_1.IN distortionUnit_2.myOpamp_0.INn VGND.t168 sky130_fd_pr__res_xhigh_po_0p35 l=10
X98 VPWR.t294 a_20584_23723# a_20584_23723# VPWR.t293 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X99 VGND.t382 VGND.t380 VGND.t381 VGND.t310 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0 ps=0 w=0.42 l=1
X100 a_20584_23723# distortionUnit_6.IN a_20842_23723# VGND.t212 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X101 a_20934_16677# distortionUnit_7.IN a_21192_16677# VGND.t61 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X102 a_20584_23723# VGND.t378 VGND.t379 VGND.t288 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X103 distortionUnit_2.tgate_1.CTRLB ui_in[1].t4 VPWR.t84 distortionUnit_2.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X104 distortionUnit_4.tgate_1.CTRLB ui_in[3].t5 VGND.t63 VGND.t62 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X105 distortionUnit_0.tgate_1.IN a_7752_16807# VPWR.t45 VPWR.t44 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X106 VGND.t416 ui_in[5].t3 distortionUnit_6.tgate_1.CTRLB VGND.t415 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X107 VPWR.t297 ui_in[6].t5 distortionUnit_0.tgate_1.CTRLB distortionUnit_0.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X108 distortionUnit_7.tgate_1.CTRLB ui_in[7].t2 VPWR.t300 distortionUnit_7.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X109 VPWR.t191 ui_in[7].t3 distortionUnit_7.tgate_1.CTRLB distortionUnit_7.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X110 distortionUnit_2.IN distortionUnit_1.tgate_1.CTRLB ua[0].t2 VGND.t203 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X111 distortionUnit_0.tgate_1.IN distortionUnit_0.tgate_1.CTRLB distortionUnit_7.IN VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X112 VGND.t377 VGND.t376 VGND.t377 VGND.t97 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X113 VGND.t375 VGND.t373 VGND.t375 VGND.t374 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X114 a_20746_30481# distortionUnit_4.myOpamp_0.INn distortionUnit_4.tgate_1.IN VGND.t99 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X115 VPWR.t109 a_7710_36445# a_7710_36445# VPWR.t108 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X116 distortionUnit_2.tgate_1.IN distortionUnit_2.myOpamp_0.INn a_20782_36601# VGND.t134 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X117 VPWR.t152 a_7756_30557# distortionUnit_3.tgate_1.IN VPWR.t151 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X118 VGND.t450 a_6866_35990# a_6866_35990# VGND.t54 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X119 distortionUnit_1.tgate_1.IN distortionUnit_1.tgate_1.CTRLB distortionUnit_2.IN VPWR.t180 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X120 VGND.t457 a_20090_16222# a_20090_16222# VGND.t433 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X121 VPWR.t11 ui_in[6].t6 distortionUnit_0.tgate_1.CTRLB distortionUnit_0.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X122 distortionUnit_3.tgate_1.CTRLB ui_in[2].t3 VPWR.t53 distortionUnit_3.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X123 a_7968_36445# ua[0].t4 a_7710_36445# VGND.t106 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X124 a_8014_30557# distortionUnit_3.myOpamp_0.INn distortionUnit_3.tgate_1.IN VGND.t79 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X125 distortionUnit_2.tgate_1.CTRLB ui_in[1].t5 VPWR.t192 distortionUnit_2.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X126 distortionUnit_2.tgate_1.IN a_20524_36601# VPWR.t210 VPWR.t209 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X127 VGND.t167 ui_in[3].t6 distortionUnit_4.tgate_1.CTRLB VGND.t166 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X128 VPWR.t26 a_19644_30026# VGND.t66 sky130_fd_pr__res_xhigh_po_0p35 l=0.16
X129 distortionUnit_6.OUT ui_in[5].t4 distortionUnit_6.tgate_1.IN VGND.t26 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X130 distortionUnit_2.tgate_1.IN a_20524_36601# VPWR.t208 VPWR.t207 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X131 a_20488_30481# a_20488_30481# VPWR.t175 VPWR.t174 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X132 a_20090_16222# a_20090_16222# VGND.t456 VGND.t58 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X133 a_19644_30026# a_19644_30026# VGND.t128 VGND.t127 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X134 a_20524_36601# distortionUnit_2.IN a_20782_36601# VGND.t143 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X135 distortionUnit_3.tgate_1.CTRLB ui_in[2].t4 VPWR.t303 distortionUnit_3.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X136 VPWR.t27 ui_in[2].t5 distortionUnit_3.tgate_1.CTRLB distortionUnit_3.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X137 a_7710_36445# VPWR.t256 VPWR.t258 VPWR.t257 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X138 VGND.t372 VGND.t371 distortionUnit_6.tgate_1.IN VGND.t275 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X139 distortionUnit_1.tgate_1.IN distortionUnit_1.myOpamp_0.INn a_7968_36445# VGND.t55 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X140 VGND.t370 VGND.t369 distortionUnit_5.tgate_1.IN VGND.t270 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X141 distortionUnit_7.tgate_1.IN distortionUnit_7.tgate_1.CTRLB ua[1].t3 VPWR.t158 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X142 VGND.t70 ui_in[3].t7 distortionUnit_4.tgate_1.CTRLB VGND.t69 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X143 distortionUnit_3.tgate_1.IN distortionUnit_3.myOpamp_0.INn a_8014_30557# VGND.t77 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X144 a_20842_23723# distortionUnit_6.myOpamp_0.INn distortionUnit_6.tgate_1.IN VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X145 VPWR.t70 a_7876_23853# a_7876_23853# VPWR.t69 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X146 distortionUnit_0.tgate_1.CTRLB ui_in[6].t7 VPWR.t23 distortionUnit_0.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X147 VGND.t368 VGND.t366 VGND.t368 VGND.t367 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X148 a_7710_36445# ua[0].t5 a_7968_36445# VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X149 distortionUnit_6.tgate_1.CTRLB ui_in[5].t5 VGND.t40 VGND.t39 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X150 VPWR.t121 a_20934_16677# a_20934_16677# VPWR.t120 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X151 distortionUnit_3.tgate_1.IN distortionUnit_3.myOpamp_0.INn a_8014_30557# VGND.t179 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X152 distortionUnit_1.tgate_1.IN distortionUnit_1.myOpamp_0.INn VGND.t408 sky130_fd_pr__res_xhigh_po_0p35 l=10
X153 VGND.t49 a_6908_16352# a_6908_16352# VGND.t10 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X154 VPWR.t206 a_20524_36601# a_20524_36601# VPWR.t205 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X155 a_8134_23853# distortionUnit_5.IN.t12 a_7876_23853# VGND.t108 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X156 distortionUnit_7.IN ui_in[6].t8 distortionUnit_0.tgate_1.IN VGND.t207 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X157 VPWR.t204 a_20524_36601# a_20524_36601# VPWR.t203 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X158 VPWR.t5 ui_in[0].t5 distortionUnit_1.tgate_1.CTRLB distortionUnit_1.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X159 VPWR.t173 a_20488_30481# distortionUnit_4.tgate_1.IN VPWR.t172 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X160 distortionUnit_1.tgate_1.IN a_7710_36445# VPWR.t107 VPWR.t106 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X161 distortionUnit_1.tgate_1.CTRLB ui_in[0].t6 VPWR.t159 distortionUnit_1.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X162 distortionUnit_2.IN ui_in[0].t7 distortionUnit_1.tgate_1.IN VGND.t42 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X163 a_20782_36601# distortionUnit_2.myOpamp_0.INn distortionUnit_2.tgate_1.IN VGND.t133 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X164 VGND.t365 VGND.t363 VGND.t364 VGND.t278 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0 ps=0 w=0.42 l=1
X165 distortionUnit_3.tgate_1.IN distortionUnit_3.myOpamp_0.INn VGND.t27 sky130_fd_pr__res_xhigh_po_0p35 l=10
X166 distortionUnit_4.tgate_1.IN distortionUnit_4.tgate_1.CTRLB distortionUnit_5.IN.t7 VPWR.t309 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X167 ua[1].t2 distortionUnit_7.tgate_1.CTRLB distortionUnit_7.tgate_1.IN VPWR.t157 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X168 VGND.t362 VGND.t360 distortionUnit_0.tgate_1.IN VGND.t361 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X169 VGND.t146 ui_in[2].t6 distortionUnit_3.tgate_1.CTRLB VGND.t145 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X170 VGND.t359 VGND.t358 VGND.t359 VGND.t29 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X171 a_8010_16807# distortionUnit_6.OUT a_7752_16807# VGND.t50 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X172 a_20934_16677# VPWR.t253 VPWR.t255 VPWR.t254 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X173 VPWR a_6866_35990# VGND sky130_fd_pr__res_xhigh_po_0p35 l=26.11
X174 distortionUnit_0.tgate_1.IN distortionUnit_0.myOpamp_0.INn VGND.t186 sky130_fd_pr__res_xhigh_po_0p35 l=10
X175 distortionUnit_6.tgate_1.CTRLB ui_in[5].t6 VGND.t103 VGND.t102 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X176 VGND.t84 a_6912_30102# a_8014_30557# VGND.t83 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X177 VPWR.t182 a_7032_23398# VGND.t206 sky130_fd_pr__res_xhigh_po_0p35 l=0.16
X178 VGND.t357 VGND.t356 VGND.t357 VGND.t172 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X179 VGND.t197 ui_in[5].t7 distortionUnit_6.tgate_1.CTRLB VGND.t196 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X180 distortionUnit_1.tgate_1.CTRLB ui_in[0].t8 VPWR.t52 distortionUnit_1.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X181 distortionUnit_7.tgate_1.CTRLB ui_in[7].t4 VPWR.t16 distortionUnit_7.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X182 a_20524_36601# VPWR.t250 VPWR.t252 VPWR.t251 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X183 VPWR.t50 ui_in[7].t5 distortionUnit_7.tgate_1.CTRLB distortionUnit_7.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X184 VPWR.t3 a_19680_36146# VGND.t13 sky130_fd_pr__res_xhigh_po_0p35 l=0.16
X185 distortionUnit_1.tgate_1.CTRLB ui_in[0].t9 VGND.t154 VGND.t153 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X186 VGND.t418 ui_in[0].t10 distortionUnit_1.tgate_1.CTRLB VGND.t417 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X187 distortionUnit_7.IN distortionUnit_0.tgate_1.CTRLB distortionUnit_0.tgate_1.IN VPWR.t8 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X188 distortionUnit_0.tgate_1.IN distortionUnit_0.myOpamp_0.INn a_8010_16807# VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X189 distortionUnit_5.IN.t9 distortionUnit_4.tgate_1.CTRLB distortionUnit_4.IN VGND.t461 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X190 distortionUnit_3.tgate_1.CTRLB ui_in[2].t7 VGND.t412 VGND.t411 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X191 VPWR.t43 a_7752_16807# a_7752_16807# VPWR.t42 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X192 VGND.t355 VGND.t354 VGND.t355 VGND.t267 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X193 VPWR.t7 ui_in[7].t6 distortionUnit_7.tgate_1.CTRLB distortionUnit_7.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X194 VGND.t445 a_19740_23268# a_20842_23723# VGND.t210 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X195 VPWR.t14 ui_in[3].t8 distortionUnit_4.tgate_1.CTRLB distortionUnit_4.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X196 distortionUnit_4.tgate_1.IN distortionUnit_4.myOpamp_0.INn a_20746_30481# VGND.t98 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X197 ua[1].t7 ui_in[7].t7 distortionUnit_7.tgate_1.IN VGND.t95 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X198 a_21192_16677# distortionUnit_7.IN a_20934_16677# VGND.t60 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X199 distortionUnit_3.tgate_1.CTRLB ui_in[2].t8 VGND.t113 VGND.t112 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X200 VPWR.t150 a_7756_30557# a_7756_30557# VPWR.t149 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X201 a_7752_16807# VGND.t351 VGND.t353 VGND.t352 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X202 VGND.t350 VGND.t348 VGND.t350 VGND.t349 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X203 distortionUnit_2.tgate_1.CTRLB ui_in[1].t6 VPWR.t136 distortionUnit_2.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X204 distortionUnit_0.tgate_1.CTRLB ui_in[6].t9 VGND.t18 VGND.t17 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X205 VGND.t201 ui_in[0].t11 distortionUnit_1.tgate_1.CTRLB VGND.t200 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X206 VGND.t347 VGND.t346 VGND.t347 VGND.t57 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X207 VPWR.t87 ui_in[1].t7 distortionUnit_2.tgate_1.CTRLB distortionUnit_2.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X208 a_7876_23853# distortionUnit_5.IN.t13 a_8134_23853# VGND.t157 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X209 VGND.t141 a_19680_36146# a_20782_36601# VGND.t140 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X210 VGND.t345 VGND.t344 VGND.t345 VGND.t260 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X211 VPWR.t302 ui_in[7].t8 distortionUnit_7.tgate_1.CTRLB distortionUnit_7.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X212 distortionUnit_7.tgate_1.CTRLB ui_in[7].t9 VPWR.t299 distortionUnit_7.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X213 a_20746_30481# a_19644_30026# VGND.t126 VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X214 distortionUnit_2.tgate_1.IN distortionUnit_2.tgate_1.CTRLB distortionUnit_3.IN VPWR.t132 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X215 VPWR.t41 a_7752_16807# distortionUnit_0.tgate_1.IN VPWR.t40 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X216 distortionUnit_7.tgate_1.IN ui_in[7].t10 ua[1].t6 VGND.t223 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X217 a_20842_23723# a_19740_23268# VGND.t444 VGND.t28 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X218 VPWR.t222 ui_in[4].t5 distortionUnit_5.tgate_1.CTRLB distortionUnit_5.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X219 VPWR.t82 ui_in[1].t8 distortionUnit_2.tgate_1.CTRLB distortionUnit_2.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X220 VPWR.t119 a_20934_16677# distortionUnit_7.tgate_1.IN VPWR.t118 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X221 distortionUnit_4.tgate_1.CTRLB ui_in[3].t9 VPWR.t275 distortionUnit_4.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X222 VGND.t343 VGND.t341 VGND.t342 VGND.t255 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0 ps=0 w=0.42 l=1
X223 VPWR.t0 ui_in[2].t9 distortionUnit_3.tgate_1.CTRLB distortionUnit_3.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X224 a_7756_30557# a_7756_30557# VPWR.t148 VPWR.t147 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X225 distortionUnit_6.tgate_1.IN distortionUnit_6.myOpamp_0.INn a_20842_23723# VGND.t30 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X226 VPWR.t202 a_20524_36601# distortionUnit_2.tgate_1.IN VPWR.t201 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X227 VPWR.t20 ui_in[1].t9 distortionUnit_2.tgate_1.CTRLB distortionUnit_2.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X228 a_8134_23853# distortionUnit_5.myOpamp_0.INn distortionUnit_5.tgate_1.IN VGND.t155 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X229 a_8014_30557# distortionUnit_3.IN a_7756_30557# VGND.t247 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X230 distortionUnit_3.IN distortionUnit_2.tgate_1.CTRLB distortionUnit_2.IN VGND.t188 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X231 distortionUnit_3.IN distortionUnit_2.tgate_1.CTRLB distortionUnit_2.tgate_1.IN VPWR.t131 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X232 distortionUnit_0.tgate_1.IN ui_in[6].t10 distortionUnit_7.IN VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X233 distortionUnit_7.tgate_1.CTRLB ui_in[7].t11 VGND.t120 VGND.t119 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X234 VPWR.t249 VPWR.t247 distortionUnit_1.tgate_1.IN VPWR.t248 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X235 distortionUnit_0.tgate_1.IN a_7752_16807# VPWR.t39 VPWR.t38 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X236 VPWR.t13 a_20090_16222# VGND.t35 sky130_fd_pr__res_xhigh_po_0p35 l=0.16
X237 VGND.t340 VGND.t339 VGND.t340 VGND.t170 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X238 a_20746_30481# distortionUnit_4.IN a_20488_30481# VGND.t401 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X239 VPWR.t85 ui_in[2].t10 distortionUnit_3.tgate_1.CTRLB distortionUnit_3.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X240 VPWR a_6908_16352# VGND sky130_fd_pr__res_xhigh_po_0p35 l=26.11
X241 distortionUnit_4.tgate_1.IN a_20488_30481# VPWR.t171 VPWR.t170 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X242 distortionUnit_6.tgate_1.IN a_20584_23723# VPWR.t292 VPWR.t291 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X243 distortionUnit_5.IN.t2 ui_in[3].t10 distortionUnit_4.IN VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X244 a_9638_15108# distortionUnit_0.myOpamp_0.INn VGND.t431 sky130_fd_pr__res_xhigh_po_0p35 l=4
X245 distortionUnit_7.tgate_1.IN a_20934_16677# VPWR.t117 VPWR.t116 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X246 VGND.t449 a_6866_35990# a_7968_36445# VGND.t116 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X247 VPWR.t105 a_7710_36445# a_7710_36445# VPWR.t104 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X248 VGND.t338 VGND.t337 VGND.t338 VGND.t292 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X249 VPWR.t83 a_6912_30102# VGND.t111 sky130_fd_pr__res_xhigh_po_0p35 l=0.16
X250 VGND.t426 ui_in[5].t8 distortionUnit_6.tgate_1.CTRLB VGND.t425 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X251 a_20842_23723# distortionUnit_6.IN a_20584_23723# VGND.t211 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X252 a_7032_23398# a_7032_23398# VGND.t165 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X253 distortionUnit_7.tgate_1.CTRLB ui_in[7].t12 VGND.t193 VGND.t192 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X254 distortionUnit_2.IN distortionUnit_2.tgate_1.CTRLB distortionUnit_3.IN VGND.t187 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X255 VGND.t65 ui_in[7].t13 distortionUnit_7.tgate_1.CTRLB VGND.t64 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X256 a_8010_16807# a_6908_16352# VGND.t48 VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X257 distortionUnit_1.tgate_1.CTRLB ui_in[0].t12 VPWR.t21 distortionUnit_1.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X258 a_20584_23723# a_20584_23723# VPWR.t290 VPWR.t289 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X259 distortionUnit_0.tgate_1.IN distortionUnit_0.myOpamp_0.INn a_8010_16807# VGND.t10 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X260 a_20488_30481# distortionUnit_4.IN a_20746_30481# VGND.t129 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X261 a_7968_36445# a_6866_35990# VGND.t448 VGND.t53 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X262 a_21192_16677# a_20090_16222# VGND.t455 VGND.t432 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X263 VGND.t37 ui_in[5].t9 distortionUnit_6.tgate_1.CTRLB VGND.t36 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X264 VGND.t336 VGND.t334 VGND.t336 VGND.t335 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X265 distortionUnit_3.tgate_1.CTRLB ui_in[2].t11 VGND.t110 VGND.t109 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X266 a_7968_36445# a_6866_35990# VGND.t447 VGND.t52 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X267 distortionUnit_0.tgate_1.CTRLB ui_in[6].t11 VGND.t1 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X268 VGND.t162 a_7032_23398# a_8134_23853# VGND.t161 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X269 a_7756_30557# distortionUnit_3.IN a_8014_30557# VGND.t87 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X270 a_22470_22024# distortionUnit_6.myOpamp_0.INn VGND.t407 sky130_fd_pr__res_xhigh_po_0p35 l=4
X271 a_20934_16677# distortionUnit_7.IN a_21192_16677# VGND.t59 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X272 VGND.t333 VGND.t330 VGND.t332 VGND.t331 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0 ps=0 w=0.42 l=1
X273 a_22374_28782# distortionUnit_4.myOpamp_0.INn VGND.t121 sky130_fd_pr__res_xhigh_po_0p35 l=4
X274 VPWR.t306 ui_in[0].t13 distortionUnit_1.tgate_1.CTRLB distortionUnit_1.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X275 VGND.t105 ui_in[0].t14 distortionUnit_1.tgate_1.CTRLB VGND.t104 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X276 distortionUnit_4.tgate_1.IN distortionUnit_4.myOpamp_0.INn VGND.t178 sky130_fd_pr__res_xhigh_po_0p35 l=10
X277 VPWR a_19740_23268# VGND sky130_fd_pr__res_xhigh_po_0p35 l=26.11
X278 distortionUnit_1.tgate_1.CTRLB ui_in[0].t15 VGND.t152 VGND.t151 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X279 distortionUnit_3.tgate_1.CTRLB ui_in[2].t12 VGND.t184 VGND.t183 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X280 VGND.t329 VGND.t328 VGND.t329 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X281 VPWR.t169 a_20488_30481# a_20488_30481# VPWR.t168 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X282 VGND.t177 ui_in[2].t13 distortionUnit_3.tgate_1.CTRLB VGND.t176 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X283 VGND.t125 a_19644_30026# a_19644_30026# VGND.t100 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X284 a_20782_36601# distortionUnit_2.IN a_20524_36601# VGND.t172 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X285 VPWR.t81 ui_in[3].t11 distortionUnit_4.tgate_1.CTRLB distortionUnit_4.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X286 VPWR.t288 a_20584_23723# distortionUnit_6.tgate_1.IN VPWR.t287 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X287 distortionUnit_6.IN ui_in[4].t6 distortionUnit_5.IN.t5 VPWR.t221 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X288 VGND.t218 ui_in[6].t12 distortionUnit_0.tgate_1.CTRLB VGND.t217 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X289 a_7710_36445# a_7710_36445# VPWR.t103 VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X290 distortionUnit_4.tgate_1.CTRLB ui_in[3].t12 VPWR.t188 distortionUnit_4.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X291 VGND.t327 VGND.t326 VGND.t327 VGND.t56 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X292 VGND.t325 VGND.t323 VGND.t325 VGND.t324 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X293 distortionUnit_6.tgate_1.CTRLB ui_in[5].t10 VGND.t148 VGND.t147 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X294 a_21192_16677# distortionUnit_7.myOpamp_0.INn distortionUnit_7.tgate_1.IN VGND.t434 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X295 VGND.t191 ui_in[6].t13 distortionUnit_0.tgate_1.CTRLB VGND.t190 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X296 a_7968_36445# ua[0].t6 a_7710_36445# VGND.t101 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X297 distortionUnit_1.tgate_1.CTRLB ui_in[0].t16 VGND.t429 VGND.t428 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X298 VPWR.t79 ui_in[1].t10 distortionUnit_2.tgate_1.CTRLB distortionUnit_2.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X299 a_8014_30557# distortionUnit_3.myOpamp_0.INn distortionUnit_3.tgate_1.IN VGND.t85 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X300 distortionUnit_2.tgate_1.CTRLB ui_in[1].t11 VPWR.t305 distortionUnit_2.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X301 a_8134_23853# distortionUnit_5.IN.t14 a_7876_23853# VGND.t173 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X302 distortionUnit_2.tgate_1.IN a_20524_36601# VPWR.t200 VPWR.t199 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X303 a_20488_30481# a_20488_30481# VPWR.t167 VPWR.t166 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X304 distortionUnit_5.IN.t11 distortionUnit_5.tgate_1.CTRLB distortionUnit_6.IN VGND.t463 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X305 VPWR.t101 a_7710_36445# distortionUnit_1.tgate_1.IN VPWR.t100 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X306 distortionUnit_6.tgate_1.CTRLB ui_in[5].t11 VPWR.t75 distortionUnit_6.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X307 VGND.t322 VGND.t320 VGND.t322 VGND.t321 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X308 a_20524_36601# distortionUnit_2.IN a_20782_36601# VGND.t140 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X309 distortionUnit_4.tgate_1.CTRLB ui_in[3].t13 VPWR.t130 distortionUnit_4.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X310 distortionUnit_0.tgate_1.CTRLB ui_in[6].t14 VGND.t16 VGND.t15 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X311 distortionUnit_5.tgate_1.CTRLB ui_in[4].t7 VPWR.t220 distortionUnit_5.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X312 VPWR.t99 a_7710_36445# distortionUnit_1.tgate_1.IN VPWR.t98 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X313 VGND.t317 VGND.t315 VGND.t317 VGND.t316 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X314 VGND.t319 VGND.t318 VGND.t319 VGND.t32 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X315 VGND.t314 VGND.t312 distortionUnit_7.tgate_1.IN VGND.t313 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X316 a_20934_16677# a_20934_16677# VPWR.t115 VPWR.t114 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X317 a_8134_23853# a_7032_23398# VGND.t164 VGND.t163 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X318 VPWR.t68 a_7876_23853# a_7876_23853# VPWR.t67 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X319 distortionUnit_7.tgate_1.CTRLB ui_in[7].t14 VGND.t34 VGND.t33 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X320 a_6912_30102# a_6912_30102# VGND.t82 VGND.t81 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X321 VPWR.t187 a_6866_35990# VGND.t220 sky130_fd_pr__res_xhigh_po_0p35 l=0.16
X322 a_7710_36445# VGND.t309 VGND.t311 VGND.t310 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X323 VGND.t308 VGND.t307 VGND.t308 VGND.t132 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X324 VGND.t420 ui_in[7].t15 distortionUnit_7.tgate_1.CTRLB VGND.t419 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X325 a_20524_36601# a_20524_36601# VPWR.t198 VPWR.t197 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X326 VGND.t139 a_19680_36146# a_19680_36146# VGND.t131 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X327 distortionUnit_5.tgate_1.CTRLB ui_in[4].t8 VPWR.t219 distortionUnit_5.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X328 VGND.t437 ui_in[7].t16 distortionUnit_7.tgate_1.CTRLB VGND.t436 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X329 a_9642_28858# distortionUnit_3.myOpamp_0.INn VGND.t185 sky130_fd_pr__res_xhigh_po_0p35 l=4
X330 VPWR.t218 ui_in[4].t9 distortionUnit_5.tgate_1.CTRLB distortionUnit_5.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X331 distortionUnit_1.tgate_1.IN a_7710_36445# VPWR.t97 VPWR.t96 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X332 VPWR.t37 a_7752_16807# a_7752_16807# VPWR.t36 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X333 distortionUnit_5.tgate_1.IN a_7876_23853# VPWR.t66 VPWR.t65 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X334 VPWR.t19 ui_in[5].t12 distortionUnit_6.tgate_1.CTRLB distortionUnit_6.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X335 VGND.t306 VGND.t305 VGND.t306 VGND.t180 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X336 VGND.t304 VGND.t303 VGND.t304 VGND.t214 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X337 distortionUnit_7.tgate_1.IN distortionUnit_7.myOpamp_0.INn a_21192_16677# VGND.t374 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X338 distortionUnit_4.tgate_1.IN distortionUnit_4.myOpamp_0.INn a_20746_30481# VGND.t97 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X339 distortionUnit_3.IN ui_in[2].t14 distortionUnit_4.IN VPWR.t190 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X340 VGND.t160 a_7032_23398# a_7032_23398# VGND.t159 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X341 a_7876_23853# a_7876_23853# VPWR.t64 VPWR.t63 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X342 distortionUnit_6.OUT ui_in[5].t13 distortionUnit_6.IN VPWR.t77 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X343 a_19740_23268# a_19740_23268# VGND.t443 VGND.t213 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X344 distortionUnit_6.IN distortionUnit_5.tgate_1.CTRLB distortionUnit_5.tgate_1.IN VPWR.t311 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X345 a_8010_16807# distortionUnit_6.OUT a_7752_16807# VGND.t170 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X346 distortionUnit_1.tgate_1.IN distortionUnit_1.myOpamp_0.INn a_7968_36445# VGND.t54 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X347 distortionUnit_7.tgate_1.IN distortionUnit_7.myOpamp_0.INn a_21192_16677# VGND.t433 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X348 VGND.t302 VGND.t300 VGND.t302 VGND.t301 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X349 a_7876_23853# VPWR.t244 VPWR.t246 VPWR.t245 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X350 VGND.t175 ui_in[7].t17 distortionUnit_7.tgate_1.CTRLB VGND.t174 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X351 VGND.t299 VGND.t296 VGND.t298 VGND.t297 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0 ps=0 w=0.42 l=1
X352 a_19680_36146# a_19680_36146# VGND.t138 VGND.t137 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X353 distortionUnit_7.tgate_1.CTRLB ui_in[7].t18 VGND.t6 VGND.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X354 VPWR.t196 a_20524_36601# distortionUnit_2.tgate_1.IN VPWR.t195 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X355 VGND.t295 VGND.t294 VGND.t295 VGND.t171 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X356 VGND.t293 VGND.t291 distortionUnit_2.tgate_1.IN VGND.t292 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X357 a_7752_16807# a_7752_16807# VPWR.t35 VPWR.t34 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X358 VPWR.t217 ui_in[4].t10 distortionUnit_5.tgate_1.CTRLB distortionUnit_5.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X359 VGND.t124 a_19644_30026# a_20746_30481# VGND.t123 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X360 distortionUnit_5.IN.t0 ui_in[3].t14 distortionUnit_4.tgate_1.IN VGND.t435 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X361 VGND.t236 ui_in[4].t11 distortionUnit_5.tgate_1.CTRLB VGND.t235 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X362 distortionUnit_4.tgate_1.CTRLB ui_in[3].t15 VPWR.t274 distortionUnit_4.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X363 a_7752_16807# a_7752_16807# VPWR.t33 VPWR.t32 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X364 distortionUnit_4.IN distortionUnit_3.tgate_1.CTRLB distortionUnit_3.IN VGND.t74 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X365 VPWR.t243 VPWR.t241 distortionUnit_3.tgate_1.IN VPWR.t242 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X366 distortionUnit_6.IN distortionUnit_6.tgate_1.CTRLB distortionUnit_6.OUT VGND.t410 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X367 VPWR.t276 a_6908_16352# VGND.t423 sky130_fd_pr__res_xhigh_po_0p35 l=0.16
X368 VGND.t442 a_19740_23268# a_20842_23723# VGND.t212 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X369 VGND.t225 ui_in[2].t15 distortionUnit_3.tgate_1.CTRLB VGND.t224 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X370 distortionUnit_5.tgate_1.IN ui_in[4].t12 distortionUnit_6.IN VGND.t234 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X371 distortionUnit_2.tgate_1.CTRLB ui_in[1].t12 VGND.t115 VGND.t114 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X372 a_21192_16677# distortionUnit_7.IN a_20934_16677# VGND.t58 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X373 a_8010_16807# distortionUnit_0.myOpamp_0.INn distortionUnit_0.tgate_1.IN VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X374 a_20746_30481# distortionUnit_4.IN a_20488_30481# VGND.t127 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X375 VPWR.t146 a_7756_30557# a_7756_30557# VPWR.t145 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X376 VGND.t454 a_20090_16222# a_21192_16677# VGND.t61 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X377 VGND.t24 ui_in[6].t15 distortionUnit_0.tgate_1.CTRLB VGND.t23 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X378 VGND.t290 VGND.t287 VGND.t289 VGND.t288 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0 ps=0 w=0.42 l=1
X379 distortionUnit_3.tgate_1.IN distortionUnit_3.tgate_1.CTRLB distortionUnit_4.IN VPWR.t29 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X380 a_22820_14978# distortionUnit_7.myOpamp_0.INn VGND.t7 sky130_fd_pr__res_xhigh_po_0p35 l=4
X381 distortionUnit_6.tgate_1.IN distortionUnit_6.myOpamp_0.INn VGND.t14 sky130_fd_pr__res_xhigh_po_0p35 l=10
X382 VGND.t286 VGND.t284 VGND.t285 VGND.t250 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0 ps=0 w=0.42 l=1
X383 distortionUnit_5.tgate_1.IN distortionUnit_5.myOpamp_0.INn VGND.t91 sky130_fd_pr__res_xhigh_po_0p35 l=10
X384 a_8014_30557# distortionUnit_3.IN a_7756_30557# VGND.t367 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X385 distortionUnit_1.tgate_1.CTRLB ui_in[0].t17 VGND.t94 VGND.t93 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X386 VGND.t195 ui_in[2].t16 distortionUnit_3.tgate_1.CTRLB VGND.t194 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X387 a_20746_30481# a_19644_30026# VGND.t122 VGND.t99 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X388 VPWR.t31 a_7752_16807# distortionUnit_0.tgate_1.IN VPWR.t30 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X389 VPWR a_19644_30026# VGND sky130_fd_pr__res_xhigh_po_0p35 l=26.11
X390 VGND.t283 VGND.t282 VGND.t283 VGND.t169 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X391 distortionUnit_6.tgate_1.CTRLB ui_in[5].t14 VPWR.t135 distortionUnit_6.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X392 distortionUnit_3.tgate_1.IN a_7756_30557# VPWR.t144 VPWR.t143 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X393 VGND.t216 ui_in[6].t16 distortionUnit_0.tgate_1.CTRLB VGND.t215 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X394 distortionUnit_4.tgate_1.IN a_20488_30481# VPWR.t165 VPWR.t164 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X395 VPWR.t298 ui_in[3].t16 distortionUnit_4.tgate_1.CTRLB distortionUnit_4.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X396 distortionUnit_6.tgate_1.IN a_20584_23723# VPWR.t286 VPWR.t285 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X397 distortionUnit_5.IN.t6 distortionUnit_4.tgate_1.CTRLB distortionUnit_4.tgate_1.IN VPWR.t308 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X398 distortionUnit_2.tgate_1.CTRLB ui_in[1].t13 VGND.t422 VGND.t421 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X399 VGND.t281 VGND.t280 VGND.t281 VGND.t106 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X400 VPWR.t62 a_7876_23853# distortionUnit_5.tgate_1.IN VPWR.t61 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X401 distortionUnit_0.tgate_1.IN distortionUnit_0.myOpamp_0.INn a_8010_16807# VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X402 a_20488_30481# VGND.t277 VGND.t279 VGND.t278 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X403 a_8014_30557# a_6912_30102# VGND.t80 VGND.t79 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X404 a_7756_30557# VPWR.t238 VPWR.t240 VPWR.t239 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X405 VGND.t76 ui_in[0].t18 distortionUnit_1.tgate_1.CTRLB VGND.t75 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X406 distortionUnit_6.tgate_1.IN distortionUnit_6.myOpamp_0.INn a_20842_23723# VGND.t29 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X407 VPWR a_7032_23398# VGND sky130_fd_pr__res_xhigh_po_0p35 l=26.11
X408 distortionUnit_5.tgate_1.CTRLB ui_in[4].t13 VPWR.t216 distortionUnit_5.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X409 a_7756_30557# distortionUnit_3.IN a_8014_30557# VGND.t83 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X410 distortionUnit_3.IN ui_in[1].t14 distortionUnit_2.tgate_1.IN VGND.t427 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X411 VPWR.t301 ui_in[3].t17 distortionUnit_4.tgate_1.CTRLB distortionUnit_4.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X412 VGND.t47 a_6908_16352# a_8010_16807# VGND.t46 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X413 distortionUnit_6.tgate_1.CTRLB ui_in[5].t15 VPWR.t15 distortionUnit_6.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X414 VGND.t276 VGND.t274 VGND.t276 VGND.t275 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X415 VPWR.t284 a_20584_23723# a_20584_23723# VPWR.t283 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X416 VGND.t45 a_6908_16352# a_8010_16807# VGND.t44 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X417 VPWR.t18 ui_in[5].t16 distortionUnit_6.tgate_1.CTRLB distortionUnit_6.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X418 distortionUnit_4.IN distortionUnit_4.tgate_1.CTRLB distortionUnit_5.IN.t8 VGND.t460 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X419 distortionUnit_0.tgate_1.CTRLB ui_in[6].t17 VGND.t22 VGND.t21 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X420 distortionUnit_5.tgate_1.CTRLB ui_in[4].t14 VPWR.t215 distortionUnit_5.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X421 VGND.t273 VGND.t272 VGND.t273 VGND.t55 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X422 distortionUnit_5.tgate_1.IN a_7876_23853# VPWR.t60 VPWR.t59 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X423 VPWR.t113 a_20934_16677# a_20934_16677# VPWR.t112 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X424 VGND.t271 VGND.t269 VGND.t271 VGND.t270 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X425 VPWR.t163 a_20488_30481# a_20488_30481# VPWR.t162 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X426 VGND.t78 a_6912_30102# a_6912_30102# VGND.t77 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X427 a_20842_23723# a_19740_23268# VGND.t441 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X428 VPWR.t282 a_20584_23723# a_20584_23723# VPWR.t281 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X429 VGND.t268 VGND.t266 distortionUnit_1.tgate_1.IN VGND.t267 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X430 distortionUnit_4.IN ui_in[2].t17 distortionUnit_3.IN VPWR.t189 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X431 VGND.t446 a_6866_35990# a_7968_36445# VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X432 distortionUnit_5.tgate_1.IN a_7876_23853# VPWR.t58 VPWR.t57 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X433 distortionUnit_4.IN ui_in[2].t18 distortionUnit_3.tgate_1.IN VGND.t107 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X434 a_20584_23723# distortionUnit_6.IN a_20842_23723# VGND.t210 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X435 VGND.t265 VGND.t264 VGND.t265 VGND.t179 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X436 a_20782_36601# a_19680_36146# VGND.t136 VGND.t135 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X437 VGND.t263 VGND.t262 VGND.t263 VGND.t108 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X438 distortionUnit_2.tgate_1.IN ui_in[1].t15 distortionUnit_3.IN VGND.t439 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X439 a_7968_36445# ua[0].t7 a_7710_36445# VGND.t349 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X440 a_21192_16677# distortionUnit_7.IN a_20934_16677# VGND.t57 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X441 VPWR.t214 ui_in[4].t15 distortionUnit_5.tgate_1.CTRLB distortionUnit_5.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X442 VGND.t68 ui_in[3].t18 distortionUnit_4.tgate_1.CTRLB VGND.t67 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X443 a_8010_16807# a_6908_16352# VGND.t43 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X444 distortionUnit_0.tgate_1.CTRLB ui_in[6].t18 VPWR.t183 distortionUnit_0.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X445 distortionUnit_6.IN ui_in[5].t17 distortionUnit_6.OUT VPWR.t76 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X446 VGND.t261 VGND.t259 distortionUnit_4.tgate_1.IN VGND.t260 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X447 distortionUnit_2.tgate_1.IN distortionUnit_2.myOpamp_0.INn a_20782_36601# VGND.t132 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X448 a_20584_23723# a_20584_23723# VPWR.t280 VPWR.t279 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X449 distortionUnit_5.IN.t4 ui_in[4].t16 distortionUnit_6.IN VPWR.t213 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X450 a_20746_30481# distortionUnit_4.myOpamp_0.INn distortionUnit_4.tgate_1.IN VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X451 VPWR.t95 a_7710_36445# a_7710_36445# VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X452 distortionUnit_2.tgate_1.IN distortionUnit_2.myOpamp_0.INn a_20782_36601# VGND.t131 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X453 a_20488_30481# VPWR.t235 VPWR.t237 VPWR.t236 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X454 distortionUnit_3.IN distortionUnit_3.tgate_1.CTRLB distortionUnit_4.IN VGND.t73 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X455 VPWR.t142 a_7756_30557# distortionUnit_3.tgate_1.IN VPWR.t141 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X456 a_20584_23723# VPWR.t232 VPWR.t234 VPWR.t233 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X457 a_20842_23723# distortionUnit_6.myOpamp_0.INn distortionUnit_6.tgate_1.IN VGND.t28 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X458 distortionUnit_4.IN distortionUnit_3.tgate_1.CTRLB distortionUnit_3.tgate_1.IN VPWR.t28 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X459 a_20934_16677# VGND.t254 VGND.t256 VGND.t255 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X460 distortionUnit_6.OUT distortionUnit_6.tgate_1.CTRLB distortionUnit_6.IN VGND.t409 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X461 distortionUnit_4.tgate_1.CTRLB ui_in[3].t19 VGND.t90 VGND.t89 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X462 distortionUnit_6.OUT ui_in[6].t19 distortionUnit_7.IN VPWR.t22 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X463 distortionUnit_1.tgate_1.IN a_7710_36445# VPWR.t93 VPWR.t92 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X464 distortionUnit_5.tgate_1.CTRLB ui_in[4].t17 VGND.t233 VGND.t232 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X465 distortionUnit_6.IN distortionUnit_5.tgate_1.CTRLB distortionUnit_5.IN.t10 VGND.t462 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X466 VGND.t258 VGND.t257 VGND.t258 VGND.t98 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X467 a_20782_36601# distortionUnit_2.IN a_20524_36601# VGND.t137 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X468 distortionUnit_3.tgate_1.IN a_7756_30557# VPWR.t140 VPWR.t139 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X469 VGND.t253 VGND.t252 VGND.t253 VGND.t60 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X470 distortionUnit_2.tgate_1.CTRLB ui_in[1].t16 VGND.t72 VGND.t71 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X471 a_7710_36445# a_7710_36445# VPWR.t91 VPWR.t90 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X472 VGND.t150 ui_in[1].t17 distortionUnit_2.tgate_1.CTRLB VGND.t149 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X473 a_20782_36601# distortionUnit_2.IN a_20524_36601# VGND.t171 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X474 a_22410_34902# distortionUnit_2.myOpamp_0.INn VGND.t205 sky130_fd_pr__res_xhigh_po_0p35 l=4
X475 distortionUnit_3.tgate_1.IN a_7756_30557# VPWR.t138 VPWR.t137 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X476 VGND.t158 a_7032_23398# a_8134_23853# VGND.t157 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X477 a_9596_34746# distortionUnit_1.myOpamp_0.INn VGND.t202 sky130_fd_pr__res_xhigh_po_0p35 l=4
X478 a_7710_36445# ua[0].t8 a_7968_36445# VGND.t116 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X479 distortionUnit_5.tgate_1.CTRLB ui_in[4].t18 VGND.t231 VGND.t230 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X480 VPWR.t194 a_20524_36601# a_20524_36601# VPWR.t193 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X481 VGND.t229 ui_in[4].t19 distortionUnit_5.tgate_1.CTRLB VGND.t228 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X482 a_8134_23853# distortionUnit_5.IN.t15 a_7876_23853# VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X483 distortionUnit_7.IN distortionUnit_0.tgate_1.CTRLB distortionUnit_6.OUT VGND.t19 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X484 VPWR.t231 VPWR.t229 distortionUnit_4.tgate_1.IN VPWR.t230 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X485 VPWR.t228 VPWR.t226 distortionUnit_6.tgate_1.IN VPWR.t227 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X486 VGND.t414 ui_in[1].t18 distortionUnit_2.tgate_1.CTRLB VGND.t413 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X487 VPWR.t304 ui_in[5].t18 distortionUnit_6.tgate_1.CTRLB distortionUnit_6.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X488 VPWR.t225 VPWR.t223 distortionUnit_5.tgate_1.IN VPWR.t224 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X489 VPWR.t161 a_20488_30481# distortionUnit_4.tgate_1.IN VPWR.t160 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X490 a_20524_36601# VGND.t249 VGND.t251 VGND.t250 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X491 VPWR.t278 a_20584_23723# distortionUnit_6.tgate_1.IN VPWR.t277 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X492 VPWR a_20090_16222# VGND sky130_fd_pr__res_xhigh_po_0p35 l=26.11
X493 VGND.t118 ui_in[1].t19 distortionUnit_2.tgate_1.CTRLB VGND.t117 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X494 distortionUnit_6.OUT distortionUnit_6.tgate_1.CTRLB distortionUnit_6.tgate_1.IN VPWR.t272 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X495 distortionUnit_5.tgate_1.IN distortionUnit_5.tgate_1.CTRLB distortionUnit_6.IN VPWR.t310 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X496 distortionUnit_2.IN ui_in[0].t19 ua[0].t1 VPWR.t88 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X497 distortionUnit_7.IN ui_in[7].t19 ua[1].t4 VPWR.t134 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X498 VGND.t440 a_19740_23268# a_19740_23268# VGND.t30 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X499 a_7968_36445# distortionUnit_1.myOpamp_0.INn distortionUnit_1.tgate_1.IN VGND.t53 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X500 a_21192_16677# distortionUnit_7.myOpamp_0.INn distortionUnit_7.tgate_1.IN VGND.t432 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X501 a_8010_16807# distortionUnit_6.OUT a_7752_16807# VGND.t169 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X502 distortionUnit_5.tgate_1.IN distortionUnit_5.myOpamp_0.INn a_8134_23853# VGND.t335 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X503 a_20934_16677# a_20934_16677# VPWR.t111 VPWR.t110 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X504 a_8134_23853# a_7032_23398# VGND.t156 VGND.t155 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0609 ps=0.71 w=0.42 l=1
X505 VPWR.t56 a_7876_23853# a_7876_23853# VPWR.t55 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X506 distortionUnit_3.tgate_1.IN ui_in[2].t19 distortionUnit_4.IN VGND.t38 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X507 VGND.t248 VGND.t246 VGND.t248 VGND.t247 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=1
X508 a_7968_36445# distortionUnit_1.myOpamp_0.INn distortionUnit_1.tgate_1.IN VGND.t52 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X509 VPWR.t51 ui_in[5].t19 distortionUnit_6.tgate_1.CTRLB distortionUnit_6.sky130_fd_sc_hd__tap_2_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X510 a_7876_23853# distortionUnit_5.IN.t16 a_8134_23853# VGND.t161 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X511 VPWR a_6912_30102# VGND sky130_fd_pr__res_xhigh_po_0p35 l=26.11
R0 ui_in[4].n2 ui_in[4].t9 212.081
R1 ui_in[4].n1 ui_in[4].t13 212.081
R2 ui_in[4].n6 ui_in[4].t15 212.081
R3 ui_in[4].n0 ui_in[4].t8 212.081
R4 ui_in[4].n11 ui_in[4].t10 212.081
R5 ui_in[4].n17 ui_in[4].t7 212.081
R6 ui_in[4].n12 ui_in[4].t5 212.081
R7 ui_in[4].n13 ui_in[4].t14 212.081
R8 ui_in[4] ui_in[4].n14 163.264
R9 ui_in[4].n16 ui_in[4].n15 152
R10 ui_in[4].n19 ui_in[4].n18 152
R11 ui_in[4].n10 ui_in[4].n9 152
R12 ui_in[4].n8 ui_in[4].n7 152
R13 ui_in[4].n5 ui_in[4].n4 152
R14 ui_in[4] ui_in[4].n3 152
R15 ui_in[4].n2 ui_in[4].t19 139.78
R16 ui_in[4].n1 ui_in[4].t2 139.78
R17 ui_in[4].n6 ui_in[4].t4 139.78
R18 ui_in[4].n0 ui_in[4].t18 139.78
R19 ui_in[4].n11 ui_in[4].t0 139.78
R20 ui_in[4].n17 ui_in[4].t17 139.78
R21 ui_in[4].n12 ui_in[4].t11 139.78
R22 ui_in[4].n13 ui_in[4].t3 139.78
R23 ui_in[4].n24 ui_in[4].t16 120.23
R24 ui_in[4].n24 ui_in[4].t6 120.228
R25 ui_in[4].n21 ui_in[4].t1 118.061
R26 ui_in[4].n21 ui_in[4].t12 118.058
R27 ui_in[4].n3 ui_in[4].n2 30.6732
R28 ui_in[4].n3 ui_in[4].n1 30.6732
R29 ui_in[4].n5 ui_in[4].n1 30.6732
R30 ui_in[4].n6 ui_in[4].n5 30.6732
R31 ui_in[4].n7 ui_in[4].n6 30.6732
R32 ui_in[4].n7 ui_in[4].n0 30.6732
R33 ui_in[4].n10 ui_in[4].n0 30.6732
R34 ui_in[4].n11 ui_in[4].n10 30.6732
R35 ui_in[4].n18 ui_in[4].n11 30.6732
R36 ui_in[4].n18 ui_in[4].n17 30.6732
R37 ui_in[4].n17 ui_in[4].n16 30.6732
R38 ui_in[4].n16 ui_in[4].n12 30.6732
R39 ui_in[4].n14 ui_in[4].n12 30.6732
R40 ui_in[4].n14 ui_in[4].n13 30.6732
R41 ui_in[4].n4 ui_in[4] 21.5045
R42 ui_in[4].n8 ui_in[4] 19.4565
R43 ui_in[4].n9 ui_in[4] 17.4085
R44 ui_in[4].n15 ui_in[4] 13.3125
R45 ui_in[4].n20 ui_in[4].n19 13.0565
R46 ui_in[4].n15 ui_in[4] 10.2405
R47 ui_in[4].n19 ui_in[4] 8.1925
R48 ui_in[4].n9 ui_in[4] 6.1445
R49 ui_in[4] ui_in[4].n8 4.0965
R50 ui_in[4].n23 ui_in[4].n20 3.2054
R51 ui_in[4].n20 ui_in[4] 2.3045
R52 ui_in[4].n4 ui_in[4] 2.0485
R53 ui_in[4].n22 ui_in[4].n21 0.528909
R54 ui_in[4].n25 ui_in[4].n24 0.506182
R55 ui_in[4].n26 ui_in[4].n25 0.42675
R56 ui_in[4].n26 ui_in[4].n23 0.342556
R57 ui_in[4].n23 ui_in[4].n22 0.3415
R58 ui_in[4].n25 ui_in[4] 0.170955
R59 ui_in[4].n22 ui_in[4] 0.148227
R60 ui_in[4] ui_in[4].n26 0.01225
R61 VGND.n542 VGND.n80 734302
R62 VGND.n543 VGND.n542 494301
R63 VGND.n1030 VGND.n1029 402315
R64 VGND.n1071 VGND.n52 398767
R65 VGND.n1027 VGND.n569 397435
R66 VGND.n1043 VGND.n1042 397063
R67 VGND.n265 VGND.n154 137195
R68 VGND.n366 VGND.n339 98572.6
R69 VGND.n266 VGND 82857.8
R70 VGND.n1024 VGND.n571 67471.8
R71 VGND.n1025 VGND.n569 66573.9
R72 VGND.n739 VGND.n596 54678.4
R73 VGND.n1023 VGND.n572 47151.2
R74 VGND.n157 VGND.n154 41031.3
R75 VGND.n157 VGND.n156 39882.8
R76 VGND.n234 VGND.n233 27500
R77 VGND.n486 VGND.n479 27500
R78 VGND.n724 VGND.n717 27500
R79 VGND.n807 VGND.n806 27500
R80 VGND.n997 VGND.n990 27500
R81 VGND.n944 VGND.n937 27500
R82 VGND.n308 VGND.n307 27500
R83 VGND.n431 VGND.n424 27500
R84 VGND.n841 VGND.n596 19915.8
R85 VGND.n842 VGND.n841 19476.5
R86 VGND.n1028 VGND.n1027 18975
R87 VGND.n266 VGND.n265 14154.2
R88 VGND.n234 VGND.t206 10325.8
R89 VGND.t423 VGND.n486 10325.8
R90 VGND.t220 VGND.n724 10325.8
R91 VGND.n807 VGND.t13 10325.8
R92 VGND.t111 VGND.n997 10325.8
R93 VGND.t66 VGND.n944 10325.8
R94 VGND.n308 VGND.t219 10325.8
R95 VGND.t35 VGND.n431 10325.8
R96 VGND.n246 VGND.n228 10285.8
R97 VGND.n488 VGND.n447 10285.8
R98 VGND.n726 VGND.n685 10285.8
R99 VGND.n819 VGND.n801 10285.8
R100 VGND.n999 VGND.n958 10285.8
R101 VGND.n946 VGND.n905 10285.8
R102 VGND.n320 VGND.n302 10285.8
R103 VGND.n433 VGND.n392 10285.8
R104 VGND.n235 VGND.n228 10253
R105 VGND.n485 VGND.n447 10253
R106 VGND.n723 VGND.n685 10253
R107 VGND.n808 VGND.n801 10253
R108 VGND.n996 VGND.n958 10253
R109 VGND.n943 VGND.n905 10253
R110 VGND.n309 VGND.n302 10253
R111 VGND.n430 VGND.n392 10253
R112 VGND.n246 VGND.n229 10250
R113 VGND.n488 VGND.n448 10250
R114 VGND.n726 VGND.n686 10250
R115 VGND.n819 VGND.n802 10250
R116 VGND.n999 VGND.n959 10250
R117 VGND.n946 VGND.n906 10250
R118 VGND.n320 VGND.n303 10250
R119 VGND.n433 VGND.n393 10250
R120 VGND.n235 VGND.n229 10187.3
R121 VGND.n485 VGND.n448 10187.3
R122 VGND.n723 VGND.n686 10187.3
R123 VGND.n808 VGND.n802 10187.3
R124 VGND.n996 VGND.n959 10187.3
R125 VGND.n943 VGND.n906 10187.3
R126 VGND.n309 VGND.n303 10187.3
R127 VGND.n430 VGND.n393 10187.3
R128 VGND.n565 VGND.n551 9618.24
R129 VGND.n1039 VGND.n551 9618.24
R130 VGND.n1039 VGND.n552 9618.24
R131 VGND.n546 VGND.n67 9618.24
R132 VGND.n1053 VGND.n67 9618.24
R133 VGND.n1053 VGND.n68 9618.24
R134 VGND.n164 VGND.n159 9618.24
R135 VGND.n261 VGND.n159 9618.24
R136 VGND.n261 VGND.n160 9618.24
R137 VGND.n92 VGND.n88 9618.24
R138 VGND.n534 VGND.n88 9618.24
R139 VGND.n534 VGND.n94 9618.24
R140 VGND.n606 VGND.n599 9618.24
R141 VGND.n838 VGND.n599 9618.24
R142 VGND.n838 VGND.n600 9618.24
R143 VGND.n49 VGND.n36 9618.24
R144 VGND.n1080 VGND.n36 9618.24
R145 VGND.n1080 VGND.n37 9618.24
R146 VGND.n138 VGND.n133 9618.24
R147 VGND.n335 VGND.n133 9618.24
R148 VGND.n335 VGND.n134 9618.24
R149 VGND.n372 VGND.n368 9618.24
R150 VGND.n379 VGND.n368 9618.24
R151 VGND.n379 VGND.n369 9618.24
R152 VGND.n1028 VGND.n563 9467.01
R153 VGND.n740 VGND.n739 6870.18
R154 VGND.n362 VGND.n341 6732.76
R155 VGND.n344 VGND.n343 6732.76
R156 VGND.n1066 VGND.n56 6732.76
R157 VGND.n61 VGND.n60 6732.76
R158 VGND.n767 VGND.n736 6732.76
R159 VGND.n624 VGND.n620 6732.76
R160 VGND.n1019 VGND.n575 6732.76
R161 VGND.n1013 VGND.n1008 6732.76
R162 VGND.n748 VGND.n742 6732.76
R163 VGND.n845 VGND.n583 6732.76
R164 VGND.n590 VGND.n585 6732.76
R165 VGND.n152 VGND.n146 6732.76
R166 VGND.n526 VGND.n97 6732.76
R167 VGND.n1087 VGND.n30 6732.76
R168 VGND.n544 VGND.n543 6359.87
R169 VGND.n531 VGND.n81 6141.76
R170 VGND.n540 VGND.n81 6141.76
R171 VGND.n531 VGND.n82 6141.76
R172 VGND.n540 VGND.n82 6141.76
R173 VGND.n561 VGND.n559 6141.76
R174 VGND.n1032 VGND.n559 6141.76
R175 VGND.n562 VGND.n561 6141.76
R176 VGND.n1032 VGND.n562 6141.76
R177 VGND.n77 VGND.n76 6141.76
R178 VGND.n1045 VGND.n76 6141.76
R179 VGND.n78 VGND.n77 6141.76
R180 VGND.n1045 VGND.n78 6141.76
R181 VGND.n255 VGND.n170 6141.76
R182 VGND.n255 VGND.n171 6141.76
R183 VGND.n256 VGND.n170 6141.76
R184 VGND.n256 VGND.n171 6141.76
R185 VGND.n829 VGND.n827 6141.76
R186 VGND.n831 VGND.n827 6141.76
R187 VGND.n830 VGND.n829 6141.76
R188 VGND.n831 VGND.n830 6141.76
R189 VGND.n46 VGND.n44 6141.76
R190 VGND.n1073 VGND.n44 6141.76
R191 VGND.n47 VGND.n46 6141.76
R192 VGND.n1073 VGND.n47 6141.76
R193 VGND.n329 VGND.n144 6141.76
R194 VGND.n329 VGND.n145 6141.76
R195 VGND.n330 VGND.n144 6141.76
R196 VGND.n330 VGND.n145 6141.76
R197 VGND.n131 VGND.n130 6141.76
R198 VGND.n383 VGND.n130 6141.76
R199 VGND.n382 VGND.n131 6141.76
R200 VGND.n383 VGND.n382 6141.76
R201 VGND.n563 VGND.n544 5922.05
R202 VGND.n1026 VGND.n570 5508.75
R203 VGND.n1071 VGND.n1070 5420.28
R204 VGND.n1022 VGND.n573 5159.4
R205 VGND.n1030 VGND.n563 4868.51
R206 VGND.n543 VGND.n79 4034.2
R207 VGND.n1043 VGND.n544 3806.52
R208 VGND.n1070 VGND.n53 3806.09
R209 VGND.n755 VGND.n570 3676.5
R210 VGND.n271 VGND.n270 3671.5
R211 VGND.n1069 VGND.n1068 3434.11
R212 VGND.n342 VGND.n341 3366.38
R213 VGND.n354 VGND.n343 3366.38
R214 VGND.n1066 VGND.n57 3366.38
R215 VGND.n1059 VGND.n60 3366.38
R216 VGND.n767 VGND.n737 3366.38
R217 VGND.n624 VGND.n623 3366.38
R218 VGND.n1019 VGND.n578 3366.38
R219 VGND.n1013 VGND.n1009 3366.38
R220 VGND.n748 VGND.n745 3366.38
R221 VGND.n845 VGND.n584 3366.38
R222 VGND.n590 VGND.n587 3366.38
R223 VGND.n149 VGND.n146 3366.38
R224 VGND.n526 VGND.n98 3366.38
R225 VGND.n1087 VGND.n31 3366.38
R226 VGND.n65 VGND.n54 3016.93
R227 VGND.n738 VGND 2969.99
R228 VGND.n349 VGND.n348 2399.08
R229 VGND.n594 VGND.n592 2198.58
R230 VGND.n348 VGND.n32 2191.03
R231 VGND.n1024 VGND.n1023 2145.17
R232 VGND.n270 VGND.n96 2083.37
R233 VGND.n595 VGND.n594 2036.22
R234 VGND.n751 VGND.n750 1920.23
R235 VGND.n529 VGND.n95 1850.51
R236 VGND.n366 VGND.n365 1822.86
R237 VGND.n752 VGND.n751 1776.8
R238 VGND.n756 VGND.n753 1683.19
R239 VGND.n761 VGND.n753 1683.19
R240 VGND.n616 VGND.n610 1683.19
R241 VGND.n611 VGND.n610 1683.19
R242 VGND.n1027 VGND.n1026 1503.98
R243 VGND.n1022 VGND.n1021 1499.9
R244 VGND.n351 VGND.n350 1478.96
R245 VGND.n269 VGND.n53 1460.08
R246 VGND.n1021 VGND.n574 1383.12
R247 VGND.t202 VGND.n550 1337.13
R248 VGND.n1031 VGND.t202 1337.13
R249 VGND.n351 VGND.n349 1330.05
R250 VGND.n233 VGND.t270 1302.55
R251 VGND.n479 VGND.t361 1302.55
R252 VGND.n717 VGND.t267 1302.55
R253 VGND.n806 VGND.t292 1302.55
R254 VGND.n990 VGND.t316 1302.55
R255 VGND.n937 VGND.t260 1302.55
R256 VGND.n307 VGND.t275 1302.55
R257 VGND.n424 VGND.t313 1302.55
R258 VGND.n528 VGND.n96 1281.68
R259 VGND.n592 VGND.n32 1243.6
R260 VGND.n1083 VGND.n1082 1234.1
R261 VGND.n763 VGND.n570 1234.1
R262 VGND.n1056 VGND.n1055 1234.1
R263 VGND.n1041 VGND.n549 1234.1
R264 VGND.n1028 VGND.n568 1234.1
R265 VGND.t205 VGND.n598 1231.2
R266 VGND.t205 VGND.n573 1231.2
R267 VGND.n755 VGND.n752 1229.9
R268 VGND.n750 VGND.n595 1221.82
R269 VGND.n1026 VGND.n1025 1219.12
R270 VGND.n1067 VGND.t462 1198.65
R271 VGND.n63 VGND.t463 1198.65
R272 VGND.n615 VGND.t203 1198.65
R273 VGND.t204 VGND.n612 1198.65
R274 VGND.n1020 VGND.t74 1198.65
R275 VGND.t73 VGND.n576 1198.65
R276 VGND.n749 VGND.t461 1198.65
R277 VGND.t460 VGND.n743 1198.65
R278 VGND.t188 VGND.n757 1198.65
R279 VGND.n762 VGND.t187 1198.65
R280 VGND.n591 VGND.t409 1198.65
R281 VGND.t410 VGND.n33 1198.65
R282 VGND.t19 VGND.n147 1198.65
R283 VGND.n153 VGND.t20 1198.65
R284 VGND.n346 VGND.t199 1198.65
R285 VGND.n363 VGND.t198 1198.65
R286 VGND.n263 VGND.n157 1160.48
R287 VGND.n841 VGND.n840 1083.35
R288 VGND.n337 VGND.n34 1063.33
R289 VGND.n603 VGND.n597 1063.33
R290 VGND.n264 VGND.n64 1063.33
R291 VGND.t185 VGND.n66 1055.41
R292 VGND.n1044 VGND.t185 1055.41
R293 VGND.t243 VGND.n55 1053.4
R294 VGND.t234 VGND.n1057 1053.4
R295 VGND.n766 VGND.t427 1053.4
R296 VGND.t439 VGND.n764 1053.4
R297 VGND.t42 VGND.n571 1053.4
R298 VGND.t430 VGND.n621 1053.4
R299 VGND.n1012 VGND.t107 1053.4
R300 VGND.t38 VGND.n1010 1053.4
R301 VGND.n844 VGND.t435 1053.4
R302 VGND.t189 VGND.n842 1053.4
R303 VGND.n527 VGND.t207 1053.4
R304 VGND.n156 VGND.t25 1053.4
R305 VGND.t95 VGND.n352 1053.4
R306 VGND.t223 VGND.n340 1053.4
R307 VGND.n1086 VGND.t26 1053.4
R308 VGND.t438 VGND.n1084 1053.4
R309 VGND.t121 VGND.n35 1040.9
R310 VGND.n1072 VGND.t121 1040.9
R311 VGND.t407 VGND.n132 962.694
R312 VGND.t407 VGND.n271 962.694
R313 VGND.t424 VGND.n158 962.694
R314 VGND.t424 VGND.n79 962.694
R315 VGND.n759 VGND.n753 841.596
R316 VGND.n613 VGND.n610 841.596
R317 VGND.t270 VGND.t335 803.966
R318 VGND.t335 VGND.t173 803.966
R319 VGND.t173 VGND.t157 803.966
R320 VGND.t157 VGND.t163 803.966
R321 VGND.t163 VGND.t159 803.966
R322 VGND.t2 VGND.t161 803.966
R323 VGND.t301 VGND.t155 803.966
R324 VGND.t108 VGND.t301 803.966
R325 VGND.t331 VGND.t108 803.966
R326 VGND.t361 VGND.t11 803.966
R327 VGND.t11 VGND.t169 803.966
R328 VGND.t169 VGND.t46 803.966
R329 VGND.t46 VGND.t9 803.966
R330 VGND.t9 VGND.t10 803.966
R331 VGND.t50 VGND.t44 803.966
R332 VGND.t12 VGND.t8 803.966
R333 VGND.t8 VGND.t170 803.966
R334 VGND.t170 VGND.t352 803.966
R335 VGND.t267 VGND.t55 803.966
R336 VGND.t55 VGND.t106 803.966
R337 VGND.t106 VGND.t116 803.966
R338 VGND.t116 VGND.t53 803.966
R339 VGND.t53 VGND.t54 803.966
R340 VGND.t101 VGND.t41 803.966
R341 VGND.t52 VGND.t56 803.966
R342 VGND.t56 VGND.t349 803.966
R343 VGND.t349 VGND.t310 803.966
R344 VGND.t292 VGND.t132 803.966
R345 VGND.t132 VGND.t172 803.966
R346 VGND.t172 VGND.t143 803.966
R347 VGND.t143 VGND.t135 803.966
R348 VGND.t135 VGND.t131 803.966
R349 VGND.t137 VGND.t140 803.966
R350 VGND.t134 VGND.t133 803.966
R351 VGND.t171 VGND.t134 803.966
R352 VGND.t250 VGND.t171 803.966
R353 VGND.t316 VGND.t180 803.966
R354 VGND.t180 VGND.t367 803.966
R355 VGND.t367 VGND.t87 803.966
R356 VGND.t87 VGND.t79 803.966
R357 VGND.t79 VGND.t77 803.966
R358 VGND.t81 VGND.t83 803.966
R359 VGND.t85 VGND.t179 803.966
R360 VGND.t179 VGND.t247 803.966
R361 VGND.t247 VGND.t297 803.966
R362 VGND.t260 VGND.t97 803.966
R363 VGND.t97 VGND.t401 803.966
R364 VGND.t401 VGND.t123 803.966
R365 VGND.t123 VGND.t96 803.966
R366 VGND.t96 VGND.t100 803.966
R367 VGND.t127 VGND.t129 803.966
R368 VGND.t99 VGND.t98 803.966
R369 VGND.t98 VGND.t321 803.966
R370 VGND.t321 VGND.t278 803.966
R371 VGND.t275 VGND.t32 803.966
R372 VGND.t32 VGND.t214 803.966
R373 VGND.t214 VGND.t210 803.966
R374 VGND.t210 VGND.t31 803.966
R375 VGND.t31 VGND.t30 803.966
R376 VGND.t213 VGND.t212 803.966
R377 VGND.t29 VGND.t28 803.966
R378 VGND.t211 VGND.t29 803.966
R379 VGND.t288 VGND.t211 803.966
R380 VGND.t313 VGND.t374 803.966
R381 VGND.t374 VGND.t60 803.966
R382 VGND.t60 VGND.t61 803.966
R383 VGND.t61 VGND.t432 803.966
R384 VGND.t432 VGND.t433 803.966
R385 VGND.t58 VGND.t59 803.966
R386 VGND.t434 VGND.t324 803.966
R387 VGND.t324 VGND.t57 803.966
R388 VGND.t57 VGND.t255 803.966
R389 VGND.n739 VGND.n597 795.182
R390 VGND.n542 VGND.n541 783.655
R391 VGND.n530 VGND.n529 774.306
R392 VGND.n1041 VGND 745.568
R393 VGND.n529 VGND.n528 698.878
R394 VGND.n239 VGND.n230 666.376
R395 VGND.n490 VGND.n445 666.376
R396 VGND.n728 VGND.n683 666.376
R397 VGND.n812 VGND.n803 666.376
R398 VGND.n1001 VGND.n956 666.376
R399 VGND.n948 VGND.n903 666.376
R400 VGND.n313 VGND.n304 666.376
R401 VGND.n435 VGND.n390 666.376
R402 VGND.n245 VGND.n244 665.019
R403 VGND.n489 VGND.n446 665.019
R404 VGND.n727 VGND.n684 665.019
R405 VGND.n818 VGND.n817 665.019
R406 VGND.n1000 VGND.n957 665.019
R407 VGND.n947 VGND.n904 665.019
R408 VGND.n319 VGND.n318 665.019
R409 VGND.n434 VGND.n391 665.019
R410 VGND.n238 VGND.n237 664.242
R411 VGND.n482 VGND.n480 664.242
R412 VGND.n720 VGND.n718 664.242
R413 VGND.n811 VGND.n810 664.242
R414 VGND.n993 VGND.n991 664.242
R415 VGND.n940 VGND.n938 664.242
R416 VGND.n312 VGND.n311 664.242
R417 VGND.n427 VGND.n425 664.242
R418 VGND.n236 VGND.n231 661.915
R419 VGND.n484 VGND.n483 661.915
R420 VGND.n722 VGND.n721 661.915
R421 VGND.n809 VGND.n804 661.915
R422 VGND.n995 VGND.n994 661.915
R423 VGND.n942 VGND.n941 661.915
R424 VGND.n310 VGND.n305 661.915
R425 VGND.n429 VGND.n428 661.915
R426 VGND.n268 VGND.n267 660.718
R427 VGND.t206 VGND.t331 660.674
R428 VGND.t352 VGND.t423 660.674
R429 VGND.t310 VGND.t220 660.674
R430 VGND.t13 VGND.t250 660.674
R431 VGND.t297 VGND.t111 660.674
R432 VGND.t278 VGND.t66 660.674
R433 VGND.t219 VGND.t288 660.674
R434 VGND.t255 VGND.t35 660.674
R435 VGND.n267 VGND.n53 660.265
R436 VGND.n62 VGND.t462 636.323
R437 VGND.t463 VGND.n62 636.323
R438 VGND.t203 VGND.n614 636.323
R439 VGND.n614 VGND.t204 636.323
R440 VGND.n577 VGND.t74 636.323
R441 VGND.n577 VGND.t73 636.323
R442 VGND.n744 VGND.t461 636.323
R443 VGND.n744 VGND.t460 636.323
R444 VGND.n758 VGND.t188 636.323
R445 VGND.n758 VGND.t187 636.323
R446 VGND.n586 VGND.t409 636.323
R447 VGND.n586 VGND.t410 636.323
R448 VGND.n148 VGND.t19 636.323
R449 VGND.n148 VGND.t20 636.323
R450 VGND.t199 VGND.n345 636.323
R451 VGND.n345 VGND.t198 636.323
R452 VGND.n1052 VGND.n69 632.37
R453 VGND.t161 VGND.n247 629.462
R454 VGND.n487 VGND.t44 629.462
R455 VGND.n725 VGND.t41 629.462
R456 VGND.t140 VGND.n820 629.462
R457 VGND.n998 VGND.t83 629.462
R458 VGND.n945 VGND.t129 629.462
R459 VGND.t212 VGND.n321 629.462
R460 VGND.n432 VGND.t59 629.462
R461 VGND.n260 VGND.n161 624.942
R462 VGND.n165 VGND.n161 624.942
R463 VGND.n166 VGND.n165 624.942
R464 VGND.n91 VGND.n87 624.942
R465 VGND.n91 VGND.n89 624.942
R466 VGND.n535 VGND.n87 624.942
R467 VGND.n564 VGND.n555 624.942
R468 VGND.n564 VGND.n553 624.942
R469 VGND.n1038 VGND.n553 624.942
R470 VGND.n608 VGND.n607 624.942
R471 VGND.n607 VGND.n601 624.942
R472 VGND.n837 VGND.n601 624.942
R473 VGND.n545 VGND.n73 624.942
R474 VGND.n545 VGND.n69 624.942
R475 VGND.n48 VGND.n40 624.942
R476 VGND.n48 VGND.n38 624.942
R477 VGND.n1079 VGND.n38 624.942
R478 VGND.n334 VGND.n135 624.942
R479 VGND.n139 VGND.n135 624.942
R480 VGND.n140 VGND.n139 624.942
R481 VGND.n374 VGND.n373 624.942
R482 VGND.n373 VGND.n370 624.942
R483 VGND.n378 VGND.n374 624.942
R484 VGND.n265 VGND.n264 621.763
R485 VGND.n1031 VGND.n1030 604.514
R486 VGND.n530 VGND 581.288
R487 VGND.n350 VGND 581.236
R488 VGND.n347 VGND 562.322
R489 VGND.n593 VGND 560.347
R490 VGND.n65 VGND 559.942
R491 VGND.n1058 VGND.t243 559.212
R492 VGND.n1058 VGND.t234 559.212
R493 VGND.t427 VGND.n765 559.212
R494 VGND.n765 VGND.t439 559.212
R495 VGND.n622 VGND.t42 559.212
R496 VGND.n622 VGND.t430 559.212
R497 VGND.t107 VGND.n1011 559.212
R498 VGND.n1011 VGND.t38 559.212
R499 VGND.t435 VGND.n843 559.212
R500 VGND.n843 VGND.t189 559.212
R501 VGND.n155 VGND.t207 559.212
R502 VGND.t25 VGND.n155 559.212
R503 VGND.n353 VGND.t95 559.212
R504 VGND.n353 VGND.t223 559.212
R505 VGND.t26 VGND.n1085 559.212
R506 VGND.n1085 VGND.t438 559.212
R507 VGND.n741 VGND 554.649
R508 VGND.n572 VGND 551.942
R509 VGND.n1041 VGND.n1040 529.67
R510 VGND.n1082 VGND 524.37
R511 VGND.n1055 VGND 504.416
R512 VGND.n1055 VGND.n1054 502.144
R513 VGND.n1040 VGND.n550 474.976
R514 VGND.n1082 VGND.n1081 468.348
R515 VGND.n574 VGND.n54 467.183
R516 VGND.n1072 VGND.n1071 442.577
R517 VGND.n839 VGND.n598 437.349
R518 VGND.n1044 VGND.n1043 435.115
R519 VGND.n248 VGND.t159 414.449
R520 VGND.t10 VGND.n478 414.449
R521 VGND.t54 VGND.n716 414.449
R522 VGND.n821 VGND.t131 414.449
R523 VGND.t77 VGND.n989 414.449
R524 VGND.t100 VGND.n936 414.449
R525 VGND.n322 VGND.t30 414.449
R526 VGND.t433 VGND.n423 414.449
R527 VGND.n257 VGND.n169 399.757
R528 VGND.n539 VGND.n538 399.757
R529 VGND.n1033 VGND.n558 399.757
R530 VGND.n832 VGND.n826 399.757
R531 VGND.n1046 VGND.n75 399.757
R532 VGND.n1074 VGND.n43 399.757
R533 VGND.n331 VGND.n143 399.757
R534 VGND.n384 VGND.n129 399.757
R535 VGND.n258 VGND.n257 398.683
R536 VGND.n538 VGND.n537 398.683
R537 VGND.n558 VGND.n554 398.683
R538 VGND.n826 VGND.n602 398.683
R539 VGND.n43 VGND.n39 398.683
R540 VGND.n332 VGND.n331 398.683
R541 VGND.n376 VGND.n129 398.683
R542 VGND.n248 VGND.t2 389.519
R543 VGND.n478 VGND.t50 389.519
R544 VGND.n716 VGND.t101 389.519
R545 VGND.n821 VGND.t137 389.519
R546 VGND.n989 VGND.t81 389.519
R547 VGND.n936 VGND.t127 389.519
R548 VGND.n322 VGND.t213 389.519
R549 VGND.n423 VGND.t58 389.519
R550 VGND.n1054 VGND.n66 374.904
R551 VGND.n1081 VGND.n35 369.748
R552 VGND.n1025 VGND.n1024 363.779
R553 VGND.n75 VGND.n70 349.741
R554 VGND.n572 VGND.t75 348.731
R555 VGND.n336 VGND.n132 341.969
R556 VGND.n262 VGND.n158 341.969
R557 VGND.n1023 VGND.n1022 339.307
R558 VGND.n254 VGND.n168 333.26
R559 VGND.n328 VGND.n142 333.26
R560 VGND.n375 VGND.n128 333.26
R561 VGND.n85 VGND.n84 333.26
R562 VGND.n560 VGND.n557 333.26
R563 VGND.n828 VGND.n825 333.26
R564 VGND.n45 VGND.n42 333.26
R565 VGND.n1050 VGND.n71 327.988
R566 VGND.n741 VGND.t413 319.978
R567 VGND.n259 VGND.n167 314.127
R568 VGND.n536 VGND.n86 314.127
R569 VGND.n1037 VGND.n1036 314.127
R570 VGND.n836 VGND.n835 314.127
R571 VGND.n1078 VGND.n1077 314.127
R572 VGND.n333 VGND.n141 314.127
R573 VGND.n377 VGND.n127 314.127
R574 VGND.n384 VGND.n383 292.5
R575 VGND.n383 VGND.n95 292.5
R576 VGND.n375 VGND.n131 292.5
R577 VGND.n381 VGND.n131 292.5
R578 VGND.n379 VGND.n378 292.5
R579 VGND.n380 VGND.n379 292.5
R580 VGND.n373 VGND.n372 292.5
R581 VGND.n145 VGND.n143 292.5
R582 VGND.n271 VGND.n145 292.5
R583 VGND.n144 VGND.n142 292.5
R584 VGND.n144 VGND.n132 292.5
R585 VGND.n335 VGND.n334 292.5
R586 VGND.n336 VGND.n335 292.5
R587 VGND.n139 VGND.n138 292.5
R588 VGND.n1074 VGND.n1073 292.5
R589 VGND.n1073 VGND.n1072 292.5
R590 VGND.n46 VGND.n45 292.5
R591 VGND.n46 VGND.n35 292.5
R592 VGND.n1080 VGND.n1079 292.5
R593 VGND.n1081 VGND.n1080 292.5
R594 VGND.n49 VGND.n48 292.5
R595 VGND.n832 VGND.n831 292.5
R596 VGND.n831 VGND.n573 292.5
R597 VGND.n829 VGND.n828 292.5
R598 VGND.n829 VGND.n598 292.5
R599 VGND.n838 VGND.n837 292.5
R600 VGND.n839 VGND.n838 292.5
R601 VGND.n607 VGND.n606 292.5
R602 VGND.n92 VGND.n91 292.5
R603 VGND.n171 VGND.n169 292.5
R604 VGND.n171 VGND.n79 292.5
R605 VGND.n170 VGND.n168 292.5
R606 VGND.n170 VGND.n158 292.5
R607 VGND.n261 VGND.n260 292.5
R608 VGND.n262 VGND.n261 292.5
R609 VGND.n165 VGND.n164 292.5
R610 VGND.n1046 VGND.n1045 292.5
R611 VGND.n1045 VGND.n1044 292.5
R612 VGND.n77 VGND.n72 292.5
R613 VGND.n77 VGND.n66 292.5
R614 VGND.n1053 VGND.n1052 292.5
R615 VGND.n1054 VGND.n1053 292.5
R616 VGND.n546 VGND.n545 292.5
R617 VGND.n1033 VGND.n1032 292.5
R618 VGND.n1032 VGND.n1031 292.5
R619 VGND.n561 VGND.n560 292.5
R620 VGND.n561 VGND.n550 292.5
R621 VGND.n1039 VGND.n1038 292.5
R622 VGND.n1040 VGND.n1039 292.5
R623 VGND.n565 VGND.n564 292.5
R624 VGND.n540 VGND.n539 292.5
R625 VGND.n541 VGND.n540 292.5
R626 VGND.n531 VGND.n85 292.5
R627 VGND.n532 VGND.n531 292.5
R628 VGND.n535 VGND.n534 292.5
R629 VGND.n534 VGND.n533 292.5
R630 VGND.n186 VGND.t240 287.151
R631 VGND.n115 VGND.t120 287.151
R632 VGND.n643 VGND.t154 287.151
R633 VGND.n669 VGND.t422 287.151
R634 VGND.n889 VGND.t113 287.151
R635 VGND.n863 VGND.t222 287.151
R636 VGND.n510 VGND.t18 287.151
R637 VGND.n16 VGND.t103 287.151
R638 VGND.n175 VGND.t229 284.024
R639 VGND.n104 VGND.t420 284.024
R640 VGND.n632 VGND.t76 284.024
R641 VGND.n658 VGND.t414 284.024
R642 VGND.n878 VGND.t177 284.024
R643 VGND.n852 VGND.t70 284.024
R644 VGND.n499 VGND.t218 284.024
R645 VGND.n5 VGND.t37 284.024
R646 VGND.n270 VGND.n269 278.738
R647 VGND.n372 VGND.n371 276.988
R648 VGND.n566 VGND.n565 276.257
R649 VGND.n547 VGND.n546 276.257
R650 VGND.n164 VGND.n163 276.257
R651 VGND.n93 VGND.n92 276.257
R652 VGND.n606 VGND.n605 276.257
R653 VGND.n50 VGND.n49 276.257
R654 VGND.n138 VGND.n137 276.257
R655 VGND.n840 VGND.n839 266.387
R656 VGND.t7 VGND.n381 265.567
R657 VGND.t7 VGND.n95 265.567
R658 VGND.t176 VGND.n65 265.002
R659 VGND.n1050 VGND.n1049 264.091
R660 VGND.n532 VGND.t431 263.87
R661 VGND.n541 VGND.t431 263.87
R662 VGND.n1068 VGND.n1067 261.435
R663 VGND.n1056 VGND.n63 261.435
R664 VGND.n615 VGND.n569 261.435
R665 VGND.n612 VGND.n568 261.435
R666 VGND.n1021 VGND.n1020 261.435
R667 VGND.n576 VGND.n549 261.435
R668 VGND.n750 VGND.n749 261.435
R669 VGND.n743 VGND.n596 261.435
R670 VGND.n757 VGND.n755 261.435
R671 VGND.n763 VGND.n762 261.435
R672 VGND.n592 VGND.n591 261.435
R673 VGND.n1083 VGND.n33 261.435
R674 VGND.n147 VGND.n96 261.435
R675 VGND.n154 VGND.n153 261.435
R676 VGND.n349 VGND.n346 261.435
R677 VGND.n364 VGND.n363 261.435
R678 VGND.n593 VGND.t69 260.86
R679 VGND.n137 VGND.n134 257.885
R680 VGND.n50 VGND.n37 257.885
R681 VGND.n605 VGND.n600 257.885
R682 VGND.n94 VGND.n93 257.885
R683 VGND.n163 VGND.n160 257.885
R684 VGND.n547 VGND.n68 257.885
R685 VGND.n566 VGND.n552 257.885
R686 VGND.n267 VGND 257.546
R687 VGND.n611 VGND.n609 254.685
R688 VGND.n761 VGND.n760 254.685
R689 VGND.n533 VGND 251.656
R690 VGND.n347 VGND.t36 240.785
R691 VGND.n220 VGND.t333 236.113
R692 VGND.n469 VGND.t387 236.113
R693 VGND.n707 VGND.t382 236.113
R694 VGND.n793 VGND.t286 236.113
R695 VGND.n980 VGND.t299 236.113
R696 VGND.n927 VGND.t365 236.113
R697 VGND.n294 VGND.t290 236.113
R698 VGND.n414 VGND.t343 236.113
R699 VGND.t271 VGND.n204 235.764
R700 VGND.t395 VGND.n452 235.764
R701 VGND.t355 VGND.n690 235.764
R702 VGND.t338 VGND.n777 235.764
R703 VGND.t317 VGND.n963 235.764
R704 VGND.t345 VGND.n910 235.764
R705 VGND.t276 VGND.n278 235.764
R706 VGND.t384 VGND.n397 235.764
R707 VGND.n371 VGND.n369 233.121
R708 VGND.n362 VGND.n361 232.597
R709 VGND.n355 VGND.n344 232.597
R710 VGND.n58 VGND.n56 232.597
R711 VGND.n1060 VGND.n61 232.597
R712 VGND.n736 VGND.n735 232.597
R713 VGND.n620 VGND.n619 232.597
R714 VGND.n579 VGND.n575 232.597
R715 VGND.n1008 VGND.n1007 232.597
R716 VGND.n746 VGND.n742 232.597
R717 VGND.n583 VGND.n582 232.597
R718 VGND.n588 VGND.n585 232.597
R719 VGND.n152 VGND.n151 232.597
R720 VGND.n99 VGND.n97 232.597
R721 VGND.n30 VGND.n29 232.597
R722 VGND.n1068 VGND.n55 229.755
R723 VGND.n1057 VGND.n1056 229.755
R724 VGND.n766 VGND.n752 229.755
R725 VGND.n764 VGND.n763 229.755
R726 VGND.n621 VGND.n568 229.755
R727 VGND.n1012 VGND.n574 229.755
R728 VGND.n1010 VGND.n549 229.755
R729 VGND.n844 VGND.n595 229.755
R730 VGND.n528 VGND.n527 229.755
R731 VGND.n352 VGND.n351 229.755
R732 VGND.n364 VGND.n340 229.755
R733 VGND.n1086 VGND.n32 229.755
R734 VGND.n1084 VGND.n1083 229.755
R735 VGND.n337 VGND.n336 226.944
R736 VGND.t14 VGND.n136 226.183
R737 VGND.n51 VGND.t178 226.183
R738 VGND.t168 VGND.n604 226.183
R739 VGND.t186 VGND.n90 226.183
R740 VGND.t91 VGND.n162 226.183
R741 VGND.n548 VGND.t27 226.183
R742 VGND.n567 VGND.t408 226.183
R743 VGND VGND.n339 220.334
R744 VGND.n180 VGND.n174 207.213
R745 VGND.n193 VGND.n181 207.213
R746 VGND.n183 VGND.n182 207.213
R747 VGND.n109 VGND.n103 207.213
R748 VGND.n122 VGND.n110 207.213
R749 VGND.n112 VGND.n111 207.213
R750 VGND.n637 VGND.n631 207.213
R751 VGND.n650 VGND.n638 207.213
R752 VGND.n640 VGND.n639 207.213
R753 VGND.n663 VGND.n657 207.213
R754 VGND.n676 VGND.n664 207.213
R755 VGND.n666 VGND.n665 207.213
R756 VGND.n883 VGND.n877 207.213
R757 VGND.n896 VGND.n884 207.213
R758 VGND.n886 VGND.n885 207.213
R759 VGND.n857 VGND.n851 207.213
R760 VGND.n870 VGND.n858 207.213
R761 VGND.n860 VGND.n859 207.213
R762 VGND.n504 VGND.n498 207.213
R763 VGND.n517 VGND.n505 207.213
R764 VGND.n507 VGND.n506 207.213
R765 VGND.n10 VGND.n4 207.213
R766 VGND.n23 VGND.n11 207.213
R767 VGND.n13 VGND.n12 207.213
R768 VGND.n367 VGND.n366 200.456
R769 VGND.n225 VGND.n224 194.805
R770 VGND.n474 VGND.n473 194.805
R771 VGND.n712 VGND.n711 194.805
R772 VGND.n798 VGND.n797 194.805
R773 VGND.n985 VGND.n984 194.805
R774 VGND.n932 VGND.n931 194.805
R775 VGND.n299 VGND.n298 194.805
R776 VGND.n419 VGND.n418 194.805
R777 VGND.n211 VGND.n210 194.542
R778 VGND.n459 VGND.n458 194.542
R779 VGND.n697 VGND.n696 194.542
R780 VGND.n784 VGND.n783 194.542
R781 VGND.n970 VGND.n969 194.542
R782 VGND.n917 VGND.n916 194.542
R783 VGND.n285 VGND.n284 194.542
R784 VGND.n404 VGND.n403 194.542
R785 VGND.n227 VGND.n226 194.463
R786 VGND.n213 VGND.n212 194.463
R787 VGND.n476 VGND.n475 194.463
R788 VGND.n461 VGND.n460 194.463
R789 VGND.n714 VGND.n713 194.463
R790 VGND.n699 VGND.n698 194.463
R791 VGND.n800 VGND.n799 194.463
R792 VGND.n786 VGND.n785 194.463
R793 VGND.n987 VGND.n986 194.463
R794 VGND.n972 VGND.n971 194.463
R795 VGND.n934 VGND.n933 194.463
R796 VGND.n919 VGND.n918 194.463
R797 VGND.n301 VGND.n300 194.463
R798 VGND.n287 VGND.n286 194.463
R799 VGND.n421 VGND.n420 194.463
R800 VGND.n406 VGND.n405 194.463
R801 VGND.n221 VGND.n220 194.3
R802 VGND.n223 VGND.n222 194.3
R803 VGND.n209 VGND.n208 194.3
R804 VGND.n206 VGND.n205 194.3
R805 VGND.n470 VGND.n469 194.3
R806 VGND.n472 VGND.n471 194.3
R807 VGND.n457 VGND.n456 194.3
R808 VGND.n454 VGND.n453 194.3
R809 VGND.n708 VGND.n707 194.3
R810 VGND.n710 VGND.n709 194.3
R811 VGND.n695 VGND.n694 194.3
R812 VGND.n692 VGND.n691 194.3
R813 VGND.n794 VGND.n793 194.3
R814 VGND.n796 VGND.n795 194.3
R815 VGND.n782 VGND.n781 194.3
R816 VGND.n779 VGND.n778 194.3
R817 VGND.n981 VGND.n980 194.3
R818 VGND.n983 VGND.n982 194.3
R819 VGND.n968 VGND.n967 194.3
R820 VGND.n965 VGND.n964 194.3
R821 VGND.n928 VGND.n927 194.3
R822 VGND.n930 VGND.n929 194.3
R823 VGND.n915 VGND.n914 194.3
R824 VGND.n912 VGND.n911 194.3
R825 VGND.n295 VGND.n294 194.3
R826 VGND.n297 VGND.n296 194.3
R827 VGND.n283 VGND.n282 194.3
R828 VGND.n280 VGND.n279 194.3
R829 VGND.n415 VGND.n414 194.3
R830 VGND.n417 VGND.n416 194.3
R831 VGND.n402 VGND.n401 194.3
R832 VGND.n399 VGND.n398 194.3
R833 VGND.n268 VGND.t228 190.006
R834 VGND.n233 VGND.n228 189.166
R835 VGND.n479 VGND.n447 189.166
R836 VGND.n717 VGND.n685 189.166
R837 VGND.n806 VGND.n801 189.166
R838 VGND.n990 VGND.n958 189.166
R839 VGND.n937 VGND.n905 189.166
R840 VGND.n307 VGND.n302 189.166
R841 VGND.n424 VGND.n392 189.166
R842 VGND.n338 VGND.n337 181.347
R843 VGND.n1082 VGND.n34 180.559
R844 VGND.n603 VGND.n570 180.559
R845 VGND.n1055 VGND.n64 180.559
R846 VGND.n1042 VGND.n1041 180.559
R847 VGND.n1029 VGND.n1028 180.559
R848 VGND.n247 VGND.t155 174.505
R849 VGND.n487 VGND.t12 174.505
R850 VGND.n725 VGND.t52 174.505
R851 VGND.n820 VGND.t133 174.505
R852 VGND.n998 VGND.t85 174.505
R853 VGND.n945 VGND.t99 174.505
R854 VGND.n321 VGND.t28 174.505
R855 VGND.n432 VGND.t434 174.505
R856 VGND.n594 VGND.n593 163.56
R857 VGND.n263 VGND.n262 162.695
R858 VGND.n348 VGND.n347 151.095
R859 VGND.n360 VGND.n341 147.038
R860 VGND.n1066 VGND.n1065 147.038
R861 VGND.n1061 VGND.n60 147.038
R862 VGND.n768 VGND.n767 147.038
R863 VGND.n617 VGND.n616 147.038
R864 VGND.n625 VGND.n624 147.038
R865 VGND.n1019 VGND.n1018 147.038
R866 VGND.n1014 VGND.n1013 147.038
R867 VGND.n748 VGND.n747 147.038
R868 VGND.n846 VGND.n845 147.038
R869 VGND.n756 VGND.n754 147.038
R870 VGND.n590 VGND.n589 147.038
R871 VGND.n150 VGND.n146 147.038
R872 VGND.n526 VGND.n525 147.038
R873 VGND.n356 VGND.n343 147.038
R874 VGND.n1088 VGND.n1087 147.038
R875 VGND.t75 VGND.t428 146.435
R876 VGND.t428 VGND.t200 146.435
R877 VGND.t200 VGND.t151 146.435
R878 VGND.t151 VGND.t417 146.435
R879 VGND.t417 VGND.t93 146.435
R880 VGND.n1057 VGND.n61 146.25
R881 VGND.n60 VGND.n55 146.25
R882 VGND.n63 VGND.n56 146.25
R883 VGND.n1067 VGND.n1066 146.25
R884 VGND.n764 VGND.n736 146.25
R885 VGND.n767 VGND.n766 146.25
R886 VGND.n616 VGND.n615 146.25
R887 VGND.n612 VGND.n611 146.25
R888 VGND.n621 VGND.n620 146.25
R889 VGND.n624 VGND.n571 146.25
R890 VGND.n576 VGND.n575 146.25
R891 VGND.n1020 VGND.n1019 146.25
R892 VGND.n1010 VGND.n1008 146.25
R893 VGND.n1013 VGND.n1012 146.25
R894 VGND.n743 VGND.n742 146.25
R895 VGND.n749 VGND.n748 146.25
R896 VGND.n842 VGND.n583 146.25
R897 VGND.n845 VGND.n844 146.25
R898 VGND.n757 VGND.n756 146.25
R899 VGND.n762 VGND.n761 146.25
R900 VGND.n585 VGND.n33 146.25
R901 VGND.n591 VGND.n590 146.25
R902 VGND.n153 VGND.n152 146.25
R903 VGND.n147 VGND.n146 146.25
R904 VGND.n156 VGND.n97 146.25
R905 VGND.n527 VGND.n526 146.25
R906 VGND.n344 VGND.n340 146.25
R907 VGND.n352 VGND.n343 146.25
R908 VGND.n363 VGND.n362 146.25
R909 VGND.n346 VGND.n341 146.25
R910 VGND.n1084 VGND.n30 146.25
R911 VGND.n1087 VGND.n1086 146.25
R912 VGND.t93 VGND.t104 142.615
R913 VGND.t153 VGND 141.054
R914 VGND.t413 VGND.t226 134.107
R915 VGND.t226 VGND.t149 134.107
R916 VGND.t149 VGND.t114 134.107
R917 VGND.t114 VGND.t208 134.107
R918 VGND.t208 VGND.t71 134.107
R919 VGND.t71 VGND.t117 134.107
R920 VGND.t117 VGND.n740 124.528
R921 VGND.n1069 VGND.n54 122.853
R922 VGND.n339 VGND.n338 121.493
R923 VGND.t104 VGND.t153 120.903
R924 VGND.n217 VGND.t403 118.005
R925 VGND.n203 VGND.t369 118.005
R926 VGND.n466 VGND.t351 118.005
R927 VGND.n451 VGND.t360 118.005
R928 VGND.n704 VGND.t309 118.005
R929 VGND.n689 VGND.t266 118.005
R930 VGND.n790 VGND.t249 118.005
R931 VGND.n776 VGND.t291 118.005
R932 VGND.n977 VGND.t388 118.005
R933 VGND.n962 VGND.t396 118.005
R934 VGND.n924 VGND.t277 118.005
R935 VGND.n909 VGND.t259 118.005
R936 VGND.n291 VGND.t378 118.005
R937 VGND.n277 VGND.t371 118.005
R938 VGND.n411 VGND.t254 118.005
R939 VGND.n396 VGND.t312 118.005
R940 VGND.n253 VGND.n169 111.401
R941 VGND.n327 VGND.n143 111.401
R942 VGND.n385 VGND.n384 111.401
R943 VGND.n539 VGND.n83 111.4
R944 VGND.n1034 VGND.n1033 111.4
R945 VGND.n833 VGND.n832 111.4
R946 VGND.n1047 VGND.n1046 111.4
R947 VGND.n1075 VGND.n1074 111.4
R948 VGND VGND.t112 111.335
R949 VGND.t411 VGND.t176 110.659
R950 VGND.t194 VGND.t411 110.659
R951 VGND.t183 VGND.t194 110.659
R952 VGND.t224 VGND.t183 110.659
R953 VGND.t109 VGND.t224 110.659
R954 VGND.t221 VGND 109.805
R955 VGND.t69 VGND.t62 108.898
R956 VGND.t62 VGND.t166 108.898
R957 VGND.t166 VGND.t3 108.898
R958 VGND.t3 VGND.t67 108.898
R959 VGND.t67 VGND.t89 108.898
R960 VGND.n263 VGND.n80 108.686
R961 VGND.n136 VGND.n34 108.507
R962 VGND.n52 VGND.n51 108.507
R963 VGND.n604 VGND.n603 108.507
R964 VGND.n90 VGND.n80 108.507
R965 VGND.n162 VGND.n64 108.507
R966 VGND.n1042 VGND.n548 108.507
R967 VGND.n1029 VGND.n567 108.507
R968 VGND.n260 VGND.n259 104.659
R969 VGND.n536 VGND.n535 104.659
R970 VGND.n1038 VGND.n1037 104.659
R971 VGND.n837 VGND.n836 104.659
R972 VGND.n1079 VGND.n1078 104.659
R973 VGND.n334 VGND.n333 104.659
R974 VGND.n378 VGND.n377 104.659
R975 VGND.n218 VGND.t330 104.028
R976 VGND.n216 VGND.t262 104.028
R977 VGND.n215 VGND.t300 104.028
R978 VGND.n201 VGND.t392 104.028
R979 VGND.n207 VGND.t334 104.028
R980 VGND.n202 VGND.t269 104.028
R981 VGND.n467 VGND.t385 104.028
R982 VGND.n465 VGND.t339 104.028
R983 VGND.n464 VGND.t328 104.028
R984 VGND.n449 VGND.t282 104.028
R985 VGND.n455 VGND.t390 104.028
R986 VGND.n450 VGND.t394 104.028
R987 VGND.n705 VGND.t380 104.028
R988 VGND.n703 VGND.t348 104.028
R989 VGND.n702 VGND.t326 104.028
R990 VGND.n687 VGND.t280 104.028
R991 VGND.n693 VGND.t272 104.028
R992 VGND.n688 VGND.t354 104.028
R993 VGND.n791 VGND.t284 104.028
R994 VGND.n789 VGND.t294 104.028
R995 VGND.n788 VGND.t405 104.028
R996 VGND.n774 VGND.t356 104.028
R997 VGND.n780 VGND.t307 104.028
R998 VGND.n775 VGND.t337 104.028
R999 VGND.n978 VGND.t296 104.028
R1000 VGND.n976 VGND.t246 104.028
R1001 VGND.n975 VGND.t264 104.028
R1002 VGND.n960 VGND.t366 104.028
R1003 VGND.n966 VGND.t305 104.028
R1004 VGND.n961 VGND.t315 104.028
R1005 VGND.n925 VGND.t363 104.028
R1006 VGND.n923 VGND.t320 104.028
R1007 VGND.n922 VGND.t257 104.028
R1008 VGND.n907 VGND.t400 104.028
R1009 VGND.n913 VGND.t376 104.028
R1010 VGND.n908 VGND.t344 104.028
R1011 VGND.n292 VGND.t287 104.028
R1012 VGND.n290 VGND.t398 104.028
R1013 VGND.n289 VGND.t358 104.028
R1014 VGND.n275 VGND.t303 104.028
R1015 VGND.n281 VGND.t318 104.028
R1016 VGND.n276 VGND.t274 104.028
R1017 VGND.n412 VGND.t341 104.028
R1018 VGND.n410 VGND.t346 104.028
R1019 VGND.n409 VGND.t323 104.028
R1020 VGND.n394 VGND.t252 104.028
R1021 VGND.n400 VGND.t373 104.028
R1022 VGND.n395 VGND.t383 104.028
R1023 VGND.t228 VGND.t241 100.38
R1024 VGND.t241 VGND.t237 100.38
R1025 VGND.t237 VGND.t230 100.38
R1026 VGND.t230 VGND.t244 100.38
R1027 VGND.t244 VGND.t232 100.38
R1028 VGND.t232 VGND.t235 100.38
R1029 VGND.t235 VGND.t239 100.38
R1030 VGND.t36 VGND.t147 100.38
R1031 VGND.t147 VGND.t425 100.38
R1032 VGND.t89 VGND.t181 99.3969
R1033 VGND.t239 VGND.n266 97.9907
R1034 VGND.t112 VGND.t145 95.4304
R1035 VGND.n1052 VGND.n1051 94.7205
R1036 VGND.n381 VGND.n380 94.3352
R1037 VGND.t181 VGND.t221 94.1181
R1038 VGND.n533 VGND.n532 93.7323
R1039 VGND.n751 VGND.n741 93.189
R1040 VGND.n361 VGND.n360 92.9264
R1041 VGND.n1065 VGND.n58 92.9264
R1042 VGND.n1061 VGND.n1060 92.9264
R1043 VGND.n768 VGND.n735 92.9264
R1044 VGND.n625 VGND.n619 92.9264
R1045 VGND.n1018 VGND.n579 92.9264
R1046 VGND.n1014 VGND.n1007 92.9264
R1047 VGND.n747 VGND.n746 92.9264
R1048 VGND.n846 VGND.n582 92.9264
R1049 VGND.n589 VGND.n588 92.9264
R1050 VGND.n151 VGND.n150 92.9264
R1051 VGND.n525 VGND.n99 92.9264
R1052 VGND.n356 VGND.n355 92.9264
R1053 VGND.n1088 VGND.n29 92.9264
R1054 VGND.t145 VGND.t109 92.274
R1055 VGND.n617 VGND.n609 88.4348
R1056 VGND.n760 VGND.n754 88.4348
R1057 VGND.n368 VGND.n367 87.99
R1058 VGND.n217 VGND.t404 87.6949
R1059 VGND.n466 VGND.t353 87.6949
R1060 VGND.n704 VGND.t311 87.6949
R1061 VGND.n790 VGND.t251 87.6949
R1062 VGND.n977 VGND.t389 87.6949
R1063 VGND.n924 VGND.t279 87.6949
R1064 VGND.n291 VGND.t379 87.6949
R1065 VGND.n411 VGND.t256 87.6949
R1066 VGND.n203 VGND.t370 87.5315
R1067 VGND.n451 VGND.t362 87.5315
R1068 VGND.n689 VGND.t268 87.5315
R1069 VGND.n776 VGND.t293 87.5315
R1070 VGND.n962 VGND.t397 87.5315
R1071 VGND.n909 VGND.t261 87.5315
R1072 VGND.n277 VGND.t372 87.5315
R1073 VGND.n396 VGND.t314 87.5315
R1074 VGND.t206 VGND.n229 77.0353
R1075 VGND.t423 VGND.n448 77.0353
R1076 VGND.t220 VGND.n686 77.0353
R1077 VGND.t13 VGND.n802 77.0353
R1078 VGND.t111 VGND.n959 77.0353
R1079 VGND.t66 VGND.n906 77.0353
R1080 VGND.t219 VGND.n303 77.0353
R1081 VGND.t35 VGND.n393 77.0353
R1082 VGND.t92 VGND.n338 69.1434
R1083 VGND.n167 VGND.n166 66.4099
R1084 VGND.n89 VGND.n86 66.4099
R1085 VGND.n1036 VGND.n555 66.4099
R1086 VGND.n835 VGND.n608 66.4099
R1087 VGND.n1049 VGND.n73 66.4099
R1088 VGND.n1077 VGND.n40 66.4099
R1089 VGND.n141 VGND.n140 66.4099
R1090 VGND.n370 VGND.n127 66.4099
R1091 VGND.n1059 VGND.n1058 65.0005
R1092 VGND.n62 VGND.n57 65.0005
R1093 VGND.n765 VGND.n737 65.0005
R1094 VGND.n613 VGND.n609 65.0005
R1095 VGND.n614 VGND.n613 65.0005
R1096 VGND.n623 VGND.n622 65.0005
R1097 VGND.n578 VGND.n577 65.0005
R1098 VGND.n1011 VGND.n1009 65.0005
R1099 VGND.n745 VGND.n744 65.0005
R1100 VGND.n843 VGND.n584 65.0005
R1101 VGND.n760 VGND.n759 65.0005
R1102 VGND.n759 VGND.n758 65.0005
R1103 VGND.n587 VGND.n586 65.0005
R1104 VGND.n149 VGND.n148 65.0005
R1105 VGND.n155 VGND.n98 65.0005
R1106 VGND.n354 VGND.n353 65.0005
R1107 VGND.n345 VGND.n342 65.0005
R1108 VGND.n1085 VGND.n31 65.0005
R1109 VGND.n367 VGND.n338 64.9457
R1110 VGND.n264 VGND.n263 64.2492
R1111 VGND VGND.t102 64.1195
R1112 VGND.n1060 VGND.n1059 59.3637
R1113 VGND.n58 VGND.n57 59.3637
R1114 VGND.n737 VGND.n735 59.3637
R1115 VGND.n623 VGND.n619 59.3637
R1116 VGND.n579 VGND.n578 59.3637
R1117 VGND.n1009 VGND.n1007 59.3637
R1118 VGND.n746 VGND.n745 59.3637
R1119 VGND.n584 VGND.n582 59.3637
R1120 VGND.n588 VGND.n587 59.3637
R1121 VGND.n151 VGND.n149 59.3637
R1122 VGND.n99 VGND.n98 59.3637
R1123 VGND.n355 VGND.n354 59.3637
R1124 VGND.n361 VGND.n342 59.3637
R1125 VGND.n31 VGND.n29 59.3637
R1126 VGND.n350 VGND.t419 58.4716
R1127 VGND.t217 VGND.n530 57.983
R1128 VGND.t196 VGND.t39 54.9596
R1129 VGND.t452 VGND.t196 54.9596
R1130 VGND.t415 VGND.t452 54.9596
R1131 VGND.n72 VGND.n70 49.3181
R1132 VGND.n365 VGND.t415 48.4169
R1133 VGND.n1051 VGND.n70 45.2272
R1134 VGND.n366 VGND 43.8369
R1135 VGND.n224 VGND.t156 41.4291
R1136 VGND.n224 VGND.t302 41.4291
R1137 VGND.t263 VGND.n221 41.4291
R1138 VGND.n221 VGND.t332 41.4291
R1139 VGND.t302 VGND.n223 41.4291
R1140 VGND.n223 VGND.t263 41.4291
R1141 VGND.n226 VGND.t165 41.4291
R1142 VGND.n226 VGND.t162 41.4291
R1143 VGND.n210 VGND.t393 41.4291
R1144 VGND.n210 VGND.t158 41.4291
R1145 VGND.n209 VGND.t336 41.4291
R1146 VGND.t393 VGND.n209 41.4291
R1147 VGND.n205 VGND.t271 41.4291
R1148 VGND.n205 VGND.t336 41.4291
R1149 VGND.n212 VGND.t164 41.4291
R1150 VGND.n212 VGND.t160 41.4291
R1151 VGND.n473 VGND.t43 41.4291
R1152 VGND.n473 VGND.t329 41.4291
R1153 VGND.t340 VGND.n470 41.4291
R1154 VGND.n470 VGND.t386 41.4291
R1155 VGND.t329 VGND.n472 41.4291
R1156 VGND.n472 VGND.t340 41.4291
R1157 VGND.n475 VGND.t51 41.4291
R1158 VGND.n475 VGND.t45 41.4291
R1159 VGND.n458 VGND.t283 41.4291
R1160 VGND.n458 VGND.t47 41.4291
R1161 VGND.n457 VGND.t391 41.4291
R1162 VGND.t283 VGND.n457 41.4291
R1163 VGND.n453 VGND.t395 41.4291
R1164 VGND.n453 VGND.t391 41.4291
R1165 VGND.n460 VGND.t48 41.4291
R1166 VGND.n460 VGND.t49 41.4291
R1167 VGND.n711 VGND.t447 41.4291
R1168 VGND.n711 VGND.t327 41.4291
R1169 VGND.t350 VGND.n708 41.4291
R1170 VGND.n708 VGND.t381 41.4291
R1171 VGND.t327 VGND.n710 41.4291
R1172 VGND.n710 VGND.t350 41.4291
R1173 VGND.n713 VGND.t451 41.4291
R1174 VGND.n713 VGND.t446 41.4291
R1175 VGND.n696 VGND.t281 41.4291
R1176 VGND.n696 VGND.t449 41.4291
R1177 VGND.n695 VGND.t273 41.4291
R1178 VGND.t281 VGND.n695 41.4291
R1179 VGND.n691 VGND.t355 41.4291
R1180 VGND.n691 VGND.t273 41.4291
R1181 VGND.n698 VGND.t448 41.4291
R1182 VGND.n698 VGND.t450 41.4291
R1183 VGND.n797 VGND.t142 41.4291
R1184 VGND.n797 VGND.t406 41.4291
R1185 VGND.t295 VGND.n794 41.4291
R1186 VGND.n794 VGND.t285 41.4291
R1187 VGND.t406 VGND.n796 41.4291
R1188 VGND.n796 VGND.t295 41.4291
R1189 VGND.n799 VGND.t138 41.4291
R1190 VGND.n799 VGND.t141 41.4291
R1191 VGND.n783 VGND.t357 41.4291
R1192 VGND.n783 VGND.t144 41.4291
R1193 VGND.n782 VGND.t308 41.4291
R1194 VGND.t357 VGND.n782 41.4291
R1195 VGND.n778 VGND.t338 41.4291
R1196 VGND.n778 VGND.t308 41.4291
R1197 VGND.n785 VGND.t136 41.4291
R1198 VGND.n785 VGND.t139 41.4291
R1199 VGND.n984 VGND.t86 41.4291
R1200 VGND.n984 VGND.t265 41.4291
R1201 VGND.t248 VGND.n981 41.4291
R1202 VGND.n981 VGND.t298 41.4291
R1203 VGND.t265 VGND.n983 41.4291
R1204 VGND.n983 VGND.t248 41.4291
R1205 VGND.n986 VGND.t82 41.4291
R1206 VGND.n986 VGND.t84 41.4291
R1207 VGND.n969 VGND.t368 41.4291
R1208 VGND.n969 VGND.t88 41.4291
R1209 VGND.n968 VGND.t306 41.4291
R1210 VGND.t368 VGND.n968 41.4291
R1211 VGND.n964 VGND.t317 41.4291
R1212 VGND.n964 VGND.t306 41.4291
R1213 VGND.n971 VGND.t80 41.4291
R1214 VGND.n971 VGND.t78 41.4291
R1215 VGND.n931 VGND.t122 41.4291
R1216 VGND.n931 VGND.t258 41.4291
R1217 VGND.t322 VGND.n928 41.4291
R1218 VGND.n928 VGND.t364 41.4291
R1219 VGND.t258 VGND.n930 41.4291
R1220 VGND.n930 VGND.t322 41.4291
R1221 VGND.n933 VGND.t128 41.4291
R1222 VGND.n933 VGND.t130 41.4291
R1223 VGND.n916 VGND.t402 41.4291
R1224 VGND.n916 VGND.t124 41.4291
R1225 VGND.n915 VGND.t377 41.4291
R1226 VGND.t402 VGND.n915 41.4291
R1227 VGND.n911 VGND.t345 41.4291
R1228 VGND.n911 VGND.t377 41.4291
R1229 VGND.n918 VGND.t126 41.4291
R1230 VGND.n918 VGND.t125 41.4291
R1231 VGND.n298 VGND.t444 41.4291
R1232 VGND.n298 VGND.t359 41.4291
R1233 VGND.t399 VGND.n295 41.4291
R1234 VGND.n295 VGND.t289 41.4291
R1235 VGND.t359 VGND.n297 41.4291
R1236 VGND.n297 VGND.t399 41.4291
R1237 VGND.n300 VGND.t443 41.4291
R1238 VGND.n300 VGND.t442 41.4291
R1239 VGND.n284 VGND.t304 41.4291
R1240 VGND.n284 VGND.t445 41.4291
R1241 VGND.n283 VGND.t319 41.4291
R1242 VGND.t304 VGND.n283 41.4291
R1243 VGND.n279 VGND.t276 41.4291
R1244 VGND.n279 VGND.t319 41.4291
R1245 VGND.n286 VGND.t441 41.4291
R1246 VGND.n286 VGND.t440 41.4291
R1247 VGND.n418 VGND.t458 41.4291
R1248 VGND.n418 VGND.t325 41.4291
R1249 VGND.t347 VGND.n415 41.4291
R1250 VGND.n415 VGND.t342 41.4291
R1251 VGND.t325 VGND.n417 41.4291
R1252 VGND.n417 VGND.t347 41.4291
R1253 VGND.n420 VGND.t456 41.4291
R1254 VGND.n420 VGND.t459 41.4291
R1255 VGND.n403 VGND.t253 41.4291
R1256 VGND.n403 VGND.t454 41.4291
R1257 VGND.n402 VGND.t375 41.4291
R1258 VGND.t253 VGND.n402 41.4291
R1259 VGND.n398 VGND.t384 41.4291
R1260 VGND.n398 VGND.t375 41.4291
R1261 VGND.n405 VGND.t455 41.4291
R1262 VGND.n405 VGND.t457 41.4291
R1263 VGND.t39 VGND.n364 36.6399
R1264 VGND VGND.n175 35.197
R1265 VGND VGND.n104 35.197
R1266 VGND VGND.n632 35.197
R1267 VGND VGND.n658 35.197
R1268 VGND VGND.n878 35.197
R1269 VGND VGND.n852 35.197
R1270 VGND VGND.n499 35.197
R1271 VGND VGND.n5 35.197
R1272 VGND.n179 VGND.n178 34.6358
R1273 VGND.n192 VGND.n191 34.6358
R1274 VGND.n188 VGND.n187 34.6358
R1275 VGND.n108 VGND.n107 34.6358
R1276 VGND.n121 VGND.n120 34.6358
R1277 VGND.n117 VGND.n116 34.6358
R1278 VGND.n636 VGND.n635 34.6358
R1279 VGND.n649 VGND.n648 34.6358
R1280 VGND.n645 VGND.n644 34.6358
R1281 VGND.n662 VGND.n661 34.6358
R1282 VGND.n675 VGND.n674 34.6358
R1283 VGND.n671 VGND.n670 34.6358
R1284 VGND.n882 VGND.n881 34.6358
R1285 VGND.n895 VGND.n894 34.6358
R1286 VGND.n891 VGND.n890 34.6358
R1287 VGND.n856 VGND.n855 34.6358
R1288 VGND.n869 VGND.n868 34.6358
R1289 VGND.n865 VGND.n864 34.6358
R1290 VGND.n503 VGND.n502 34.6358
R1291 VGND.n516 VGND.n515 34.6358
R1292 VGND.n512 VGND.n511 34.6358
R1293 VGND.n9 VGND.n8 34.6358
R1294 VGND.n22 VGND.n21 34.6358
R1295 VGND.n18 VGND.n17 34.6358
R1296 VGND.n254 VGND.n253 34.2005
R1297 VGND.n84 VGND.n83 34.2005
R1298 VGND.n1034 VGND.n557 34.2005
R1299 VGND.n833 VGND.n825 34.2005
R1300 VGND.n1047 VGND.n71 34.2005
R1301 VGND.n1075 VGND.n42 34.2005
R1302 VGND.n328 VGND.n327 34.2005
R1303 VGND.n385 VGND.n128 34.2005
R1304 VGND.n364 VGND.t425 33.4606
R1305 VGND.n194 VGND.n193 32.0005
R1306 VGND.n123 VGND.n122 32.0005
R1307 VGND.n651 VGND.n650 32.0005
R1308 VGND.n677 VGND.n676 32.0005
R1309 VGND.n897 VGND.n896 32.0005
R1310 VGND.n871 VGND.n870 32.0005
R1311 VGND.n518 VGND.n517 32.0005
R1312 VGND.n24 VGND.n23 32.0005
R1313 VGND.n840 VGND.n52 31.5543
R1314 VGND.n194 VGND.n180 31.2476
R1315 VGND.n123 VGND.n109 31.2476
R1316 VGND.n651 VGND.n637 31.2476
R1317 VGND.n677 VGND.n663 31.2476
R1318 VGND.n897 VGND.n883 31.2476
R1319 VGND.n871 VGND.n857 31.2476
R1320 VGND.n518 VGND.n504 31.2476
R1321 VGND.n24 VGND.n10 31.2476
R1322 VGND.t119 VGND 28.0716
R1323 VGND VGND.t17 27.836
R1324 VGND.n249 VGND.n248 26.2219
R1325 VGND.n478 VGND.n477 26.2219
R1326 VGND.n716 VGND.n715 26.2219
R1327 VGND.n822 VGND.n821 26.2219
R1328 VGND.n989 VGND.n988 26.2219
R1329 VGND.n936 VGND.n935 26.2219
R1330 VGND.n323 VGND.n322 26.2219
R1331 VGND.n423 VGND.n422 26.2219
R1332 VGND.n191 VGND.n183 25.977
R1333 VGND.n120 VGND.n112 25.977
R1334 VGND.n648 VGND.n640 25.977
R1335 VGND.n674 VGND.n666 25.977
R1336 VGND.n894 VGND.n886 25.977
R1337 VGND.n868 VGND.n860 25.977
R1338 VGND.n515 VGND.n507 25.977
R1339 VGND.n21 VGND.n13 25.977
R1340 VGND.n269 VGND.n268 25.0956
R1341 VGND.n174 VGND.t242 24.9236
R1342 VGND.n174 VGND.t238 24.9236
R1343 VGND.n181 VGND.t231 24.9236
R1344 VGND.n181 VGND.t245 24.9236
R1345 VGND.n182 VGND.t233 24.9236
R1346 VGND.n182 VGND.t236 24.9236
R1347 VGND.n103 VGND.t6 24.9236
R1348 VGND.n103 VGND.t65 24.9236
R1349 VGND.n110 VGND.t34 24.9236
R1350 VGND.n110 VGND.t175 24.9236
R1351 VGND.n111 VGND.t193 24.9236
R1352 VGND.n111 VGND.t437 24.9236
R1353 VGND.n631 VGND.t429 24.9236
R1354 VGND.n631 VGND.t201 24.9236
R1355 VGND.n638 VGND.t152 24.9236
R1356 VGND.n638 VGND.t418 24.9236
R1357 VGND.n639 VGND.t94 24.9236
R1358 VGND.n639 VGND.t105 24.9236
R1359 VGND.n657 VGND.t227 24.9236
R1360 VGND.n657 VGND.t150 24.9236
R1361 VGND.n664 VGND.t115 24.9236
R1362 VGND.n664 VGND.t209 24.9236
R1363 VGND.n665 VGND.t72 24.9236
R1364 VGND.n665 VGND.t118 24.9236
R1365 VGND.n877 VGND.t412 24.9236
R1366 VGND.n877 VGND.t195 24.9236
R1367 VGND.n884 VGND.t184 24.9236
R1368 VGND.n884 VGND.t225 24.9236
R1369 VGND.n885 VGND.t110 24.9236
R1370 VGND.n885 VGND.t146 24.9236
R1371 VGND.n851 VGND.t63 24.9236
R1372 VGND.n851 VGND.t167 24.9236
R1373 VGND.n858 VGND.t4 24.9236
R1374 VGND.n858 VGND.t68 24.9236
R1375 VGND.n859 VGND.t90 24.9236
R1376 VGND.n859 VGND.t182 24.9236
R1377 VGND.n498 VGND.t16 24.9236
R1378 VGND.n498 VGND.t216 24.9236
R1379 VGND.n505 VGND.t22 24.9236
R1380 VGND.n505 VGND.t24 24.9236
R1381 VGND.n506 VGND.t1 24.9236
R1382 VGND.n506 VGND.t191 24.9236
R1383 VGND.n4 VGND.t148 24.9236
R1384 VGND.n4 VGND.t426 24.9236
R1385 VGND.n11 VGND.t40 24.9236
R1386 VGND.n11 VGND.t197 24.9236
R1387 VGND.n12 VGND.t453 24.9236
R1388 VGND.n12 VGND.t416 24.9236
R1389 VGND.n136 VGND.n133 24.3887
R1390 VGND.n51 VGND.n36 24.3887
R1391 VGND.n604 VGND.n599 24.3887
R1392 VGND.n90 VGND.n88 24.3887
R1393 VGND.n162 VGND.n159 24.3887
R1394 VGND.n548 VGND.n67 24.3887
R1395 VGND.n567 VGND.n551 24.3887
R1396 VGND.t419 VGND.t5 24.0614
R1397 VGND.t5 VGND.t64 24.0614
R1398 VGND.t64 VGND.t33 24.0614
R1399 VGND.t33 VGND.t174 24.0614
R1400 VGND.t174 VGND.t192 24.0614
R1401 VGND.t192 VGND.t436 24.0614
R1402 VGND.t436 VGND.t119 24.0614
R1403 VGND.t15 VGND.t217 23.8595
R1404 VGND.t215 VGND.t15 23.8595
R1405 VGND.t21 VGND.t215 23.8595
R1406 VGND.t23 VGND.t21 23.8595
R1407 VGND.t0 VGND.t23 23.8595
R1408 VGND.t190 VGND.t0 23.8595
R1409 VGND.t17 VGND.t190 23.8595
R1410 VGND.n840 VGND.n597 23.8559
R1411 VGND.n382 VGND.n129 23.4005
R1412 VGND.n382 VGND.t7 23.4005
R1413 VGND.n130 VGND.n128 23.4005
R1414 VGND.t7 VGND.n130 23.4005
R1415 VGND.n331 VGND.n330 23.4005
R1416 VGND.n330 VGND.t407 23.4005
R1417 VGND.n329 VGND.n328 23.4005
R1418 VGND.t407 VGND.n329 23.4005
R1419 VGND.n47 VGND.n43 23.4005
R1420 VGND.t121 VGND.n47 23.4005
R1421 VGND.n44 VGND.n42 23.4005
R1422 VGND.t121 VGND.n44 23.4005
R1423 VGND.n830 VGND.n826 23.4005
R1424 VGND.n830 VGND.t205 23.4005
R1425 VGND.n827 VGND.n825 23.4005
R1426 VGND.t205 VGND.n827 23.4005
R1427 VGND.n257 VGND.n256 23.4005
R1428 VGND.n256 VGND.t424 23.4005
R1429 VGND.n255 VGND.n254 23.4005
R1430 VGND.t424 VGND.n255 23.4005
R1431 VGND.n78 VGND.n75 23.4005
R1432 VGND.t185 VGND.n78 23.4005
R1433 VGND.n76 VGND.n71 23.4005
R1434 VGND.t185 VGND.n76 23.4005
R1435 VGND.n562 VGND.n558 23.4005
R1436 VGND.t202 VGND.n562 23.4005
R1437 VGND.n559 VGND.n557 23.4005
R1438 VGND.t202 VGND.n559 23.4005
R1439 VGND.n538 VGND.n82 23.4005
R1440 VGND.n82 VGND.t431 23.4005
R1441 VGND.n84 VGND.n81 23.4005
R1442 VGND.n81 VGND.t431 23.4005
R1443 VGND.n231 VGND.n229 20.8934
R1444 VGND.n238 VGND.n228 20.8934
R1445 VGND.n483 VGND.n448 20.8934
R1446 VGND.n480 VGND.n447 20.8934
R1447 VGND.n721 VGND.n686 20.8934
R1448 VGND.n718 VGND.n685 20.8934
R1449 VGND.n804 VGND.n802 20.8934
R1450 VGND.n811 VGND.n801 20.8934
R1451 VGND.n994 VGND.n959 20.8934
R1452 VGND.n991 VGND.n958 20.8934
R1453 VGND.n941 VGND.n906 20.8934
R1454 VGND.n938 VGND.n905 20.8934
R1455 VGND.n305 VGND.n303 20.8934
R1456 VGND.n312 VGND.n302 20.8934
R1457 VGND.n428 VGND.n393 20.8934
R1458 VGND.n425 VGND.n392 20.8934
R1459 VGND.n266 VGND 19.1205
R1460 VGND.n178 VGND.n175 18.824
R1461 VGND.n107 VGND.n104 18.824
R1462 VGND.n635 VGND.n632 18.824
R1463 VGND.n661 VGND.n658 18.824
R1464 VGND.n881 VGND.n878 18.824
R1465 VGND.n855 VGND.n852 18.824
R1466 VGND.n502 VGND.n499 18.824
R1467 VGND.n8 VGND.n5 18.824
R1468 VGND.n370 VGND.n369 13.6052
R1469 VGND.n374 VGND.n368 13.6052
R1470 VGND.n140 VGND.n134 13.6052
R1471 VGND.n135 VGND.n133 13.6052
R1472 VGND.n40 VGND.n37 13.6052
R1473 VGND.n38 VGND.n36 13.6052
R1474 VGND.n608 VGND.n600 13.6052
R1475 VGND.n601 VGND.n599 13.6052
R1476 VGND.n94 VGND.n89 13.6052
R1477 VGND.n88 VGND.n87 13.6052
R1478 VGND.n166 VGND.n160 13.6052
R1479 VGND.n161 VGND.n159 13.6052
R1480 VGND.n73 VGND.n68 13.6052
R1481 VGND.n69 VGND.n67 13.6052
R1482 VGND.n555 VGND.n552 13.6052
R1483 VGND.n553 VGND.n551 13.6052
R1484 VGND.n187 VGND.n186 13.5534
R1485 VGND.n116 VGND.n115 13.5534
R1486 VGND.n644 VGND.n643 13.5534
R1487 VGND.n670 VGND.n669 13.5534
R1488 VGND.n890 VGND.n889 13.5534
R1489 VGND.n864 VGND.n863 13.5534
R1490 VGND.n511 VGND.n510 13.5534
R1491 VGND.n17 VGND.n16 13.5534
R1492 VGND.n380 VGND.n338 12.5785
R1493 VGND.n360 VGND 11.4981
R1494 VGND.n1065 VGND 11.4981
R1495 VGND VGND.n1061 11.4981
R1496 VGND VGND.n768 11.4981
R1497 VGND VGND.n617 11.4981
R1498 VGND VGND.n625 11.4981
R1499 VGND.n1018 VGND 11.4981
R1500 VGND VGND.n1014 11.4981
R1501 VGND.n747 VGND 11.4981
R1502 VGND VGND.n846 11.4981
R1503 VGND.n754 VGND 11.4981
R1504 VGND.n589 VGND 11.4981
R1505 VGND.n150 VGND 11.4981
R1506 VGND.n525 VGND 11.4981
R1507 VGND VGND.n356 11.4981
R1508 VGND VGND.n1088 11.4981
R1509 VGND.n186 VGND.n185 11.1829
R1510 VGND.n115 VGND.n114 11.1829
R1511 VGND.n643 VGND.n642 11.1829
R1512 VGND.n669 VGND.n668 11.1829
R1513 VGND.n889 VGND.n888 11.1829
R1514 VGND.n863 VGND.n862 11.1829
R1515 VGND.n510 VGND.n509 11.1829
R1516 VGND.n16 VGND.n15 11.1829
R1517 VGND.n1070 VGND.n1069 11.1086
R1518 VGND.n1051 VGND.n1050 10.1983
R1519 VGND.n176 VGND.n175 9.3005
R1520 VGND.n178 VGND.n177 9.3005
R1521 VGND.n179 VGND.n172 9.3005
R1522 VGND.n195 VGND.n194 9.3005
R1523 VGND.n192 VGND.n173 9.3005
R1524 VGND.n191 VGND.n190 9.3005
R1525 VGND.n189 VGND.n188 9.3005
R1526 VGND.n187 VGND.n184 9.3005
R1527 VGND.n105 VGND.n104 9.3005
R1528 VGND.n107 VGND.n106 9.3005
R1529 VGND.n108 VGND.n101 9.3005
R1530 VGND.n124 VGND.n123 9.3005
R1531 VGND.n121 VGND.n102 9.3005
R1532 VGND.n120 VGND.n119 9.3005
R1533 VGND.n118 VGND.n117 9.3005
R1534 VGND.n116 VGND.n113 9.3005
R1535 VGND.n633 VGND.n632 9.3005
R1536 VGND.n635 VGND.n634 9.3005
R1537 VGND.n636 VGND.n629 9.3005
R1538 VGND.n652 VGND.n651 9.3005
R1539 VGND.n649 VGND.n630 9.3005
R1540 VGND.n648 VGND.n647 9.3005
R1541 VGND.n646 VGND.n645 9.3005
R1542 VGND.n644 VGND.n641 9.3005
R1543 VGND.n659 VGND.n658 9.3005
R1544 VGND.n661 VGND.n660 9.3005
R1545 VGND.n662 VGND.n655 9.3005
R1546 VGND.n678 VGND.n677 9.3005
R1547 VGND.n675 VGND.n656 9.3005
R1548 VGND.n674 VGND.n673 9.3005
R1549 VGND.n672 VGND.n671 9.3005
R1550 VGND.n670 VGND.n667 9.3005
R1551 VGND.n879 VGND.n878 9.3005
R1552 VGND.n881 VGND.n880 9.3005
R1553 VGND.n882 VGND.n875 9.3005
R1554 VGND.n898 VGND.n897 9.3005
R1555 VGND.n895 VGND.n876 9.3005
R1556 VGND.n894 VGND.n893 9.3005
R1557 VGND.n892 VGND.n891 9.3005
R1558 VGND.n890 VGND.n887 9.3005
R1559 VGND.n853 VGND.n852 9.3005
R1560 VGND.n855 VGND.n854 9.3005
R1561 VGND.n856 VGND.n849 9.3005
R1562 VGND.n872 VGND.n871 9.3005
R1563 VGND.n869 VGND.n850 9.3005
R1564 VGND.n868 VGND.n867 9.3005
R1565 VGND.n866 VGND.n865 9.3005
R1566 VGND.n864 VGND.n861 9.3005
R1567 VGND.n500 VGND.n499 9.3005
R1568 VGND.n502 VGND.n501 9.3005
R1569 VGND.n503 VGND.n496 9.3005
R1570 VGND.n519 VGND.n518 9.3005
R1571 VGND.n516 VGND.n497 9.3005
R1572 VGND.n515 VGND.n514 9.3005
R1573 VGND.n513 VGND.n512 9.3005
R1574 VGND.n511 VGND.n508 9.3005
R1575 VGND.n6 VGND.n5 9.3005
R1576 VGND.n8 VGND.n7 9.3005
R1577 VGND.n9 VGND.n2 9.3005
R1578 VGND.n25 VGND.n24 9.3005
R1579 VGND.n22 VGND.n3 9.3005
R1580 VGND.n21 VGND.n20 9.3005
R1581 VGND.n19 VGND.n18 9.3005
R1582 VGND.n17 VGND.n14 9.3005
R1583 VGND.n188 VGND.n183 8.65932
R1584 VGND.n117 VGND.n112 8.65932
R1585 VGND.n645 VGND.n640 8.65932
R1586 VGND.n671 VGND.n666 8.65932
R1587 VGND.n891 VGND.n886 8.65932
R1588 VGND.n865 VGND.n860 8.65932
R1589 VGND.n512 VGND.n507 8.65932
R1590 VGND.n18 VGND.n13 8.65932
R1591 VGND.n740 VGND.n738 8.57205
R1592 VGND.n236 VGND.n235 8.23994
R1593 VGND.n235 VGND.n234 8.23994
R1594 VGND.n246 VGND.n245 8.23994
R1595 VGND.n247 VGND.n246 8.23994
R1596 VGND.n485 VGND.n484 8.23994
R1597 VGND.n486 VGND.n485 8.23994
R1598 VGND.n489 VGND.n488 8.23994
R1599 VGND.n488 VGND.n487 8.23994
R1600 VGND.n723 VGND.n722 8.23994
R1601 VGND.n724 VGND.n723 8.23994
R1602 VGND.n727 VGND.n726 8.23994
R1603 VGND.n726 VGND.n725 8.23994
R1604 VGND.n809 VGND.n808 8.23994
R1605 VGND.n808 VGND.n807 8.23994
R1606 VGND.n819 VGND.n818 8.23994
R1607 VGND.n820 VGND.n819 8.23994
R1608 VGND.n996 VGND.n995 8.23994
R1609 VGND.n997 VGND.n996 8.23994
R1610 VGND.n1000 VGND.n999 8.23994
R1611 VGND.n999 VGND.n998 8.23994
R1612 VGND.n943 VGND.n942 8.23994
R1613 VGND.n944 VGND.n943 8.23994
R1614 VGND.n947 VGND.n946 8.23994
R1615 VGND.n946 VGND.n945 8.23994
R1616 VGND.n310 VGND.n309 8.23994
R1617 VGND.n309 VGND.n308 8.23994
R1618 VGND.n320 VGND.n319 8.23994
R1619 VGND.n321 VGND.n320 8.23994
R1620 VGND.n430 VGND.n429 8.23994
R1621 VGND.n431 VGND.n430 8.23994
R1622 VGND.n434 VGND.n433 8.23994
R1623 VGND.n433 VGND.n432 8.23994
R1624 VGND.n137 VGND.t14 7.84349
R1625 VGND.t178 VGND.n50 7.84349
R1626 VGND.n605 VGND.t168 7.84349
R1627 VGND.n93 VGND.t186 7.84349
R1628 VGND.n163 VGND.t91 7.84349
R1629 VGND.t27 VGND.n547 7.84349
R1630 VGND.t408 VGND.n566 7.84349
R1631 VGND.n371 VGND.t92 7.09041
R1632 VGND.t102 VGND.n365 6.54325
R1633 VGND.n259 VGND.n258 5.9205
R1634 VGND.n537 VGND.n536 5.9205
R1635 VGND.n1037 VGND.n554 5.9205
R1636 VGND.n836 VGND.n602 5.9205
R1637 VGND.n1078 VGND.n39 5.9205
R1638 VGND.n333 VGND.n332 5.9205
R1639 VGND.n377 VGND.n376 5.9205
R1640 VGND.n771 VGND 5.54759
R1641 VGND.n1050 VGND.n72 5.27109
R1642 VGND.n580 VGND 4.6065
R1643 VGND.n1092 VGND 3.54117
R1644 VGND.n770 VGND.n734 3.45067
R1645 VGND.n359 VGND.n358 3.45067
R1646 VGND.n1064 VGND.n1063 3.45067
R1647 VGND.n627 VGND.n618 3.45067
R1648 VGND.n1017 VGND.n1016 3.45067
R1649 VGND.n848 VGND.n581 3.45067
R1650 VGND.n523 VGND.n100 3.45067
R1651 VGND.n1090 VGND.n28 3.45067
R1652 VGND.n180 VGND.n179 3.38874
R1653 VGND.n109 VGND.n108 3.38874
R1654 VGND.n637 VGND.n636 3.38874
R1655 VGND.n663 VGND.n662 3.38874
R1656 VGND.n883 VGND.n882 3.38874
R1657 VGND.n857 VGND.n856 3.38874
R1658 VGND.n504 VGND.n503 3.38874
R1659 VGND.n10 VGND.n9 3.38874
R1660 VGND.n1063 VGND.n1062 2.87883
R1661 VGND.n770 VGND.n769 2.87883
R1662 VGND.n627 VGND.n626 2.87883
R1663 VGND.n1016 VGND.n1015 2.87883
R1664 VGND.n848 VGND.n847 2.87883
R1665 VGND.n524 VGND.n523 2.87883
R1666 VGND.n358 VGND.n357 2.87883
R1667 VGND.n1090 VGND.n1089 2.87883
R1668 VGND.n193 VGND.n192 2.63579
R1669 VGND.n122 VGND.n121 2.63579
R1670 VGND.n650 VGND.n649 2.63579
R1671 VGND.n676 VGND.n675 2.63579
R1672 VGND.n896 VGND.n895 2.63579
R1673 VGND.n870 VGND.n869 2.63579
R1674 VGND.n517 VGND.n516 2.63579
R1675 VGND.n23 VGND.n22 2.63579
R1676 VGND.n1093 VGND 2.47583
R1677 VGND.n252 VGND.n167 2.45057
R1678 VGND.n441 VGND.n86 2.45057
R1679 VGND.n1036 VGND.n1035 2.45057
R1680 VGND.n835 VGND.n834 2.45057
R1681 VGND.n1049 VGND.n1048 2.45057
R1682 VGND.n1077 VGND.n1076 2.45057
R1683 VGND.n326 VGND.n141 2.45057
R1684 VGND.n386 VGND.n127 2.45057
R1685 VGND.n1095 VGND 2.2565
R1686 VGND.n243 VGND.n232 2.09737
R1687 VGND.n243 VGND.n242 2.09737
R1688 VGND.n481 VGND.n444 2.09737
R1689 VGND.n491 VGND.n444 2.09737
R1690 VGND.n719 VGND.n682 2.09737
R1691 VGND.n729 VGND.n682 2.09737
R1692 VGND.n816 VGND.n805 2.09737
R1693 VGND.n816 VGND.n815 2.09737
R1694 VGND.n992 VGND.n955 2.09737
R1695 VGND.n1002 VGND.n955 2.09737
R1696 VGND.n939 VGND.n902 2.09737
R1697 VGND.n949 VGND.n902 2.09737
R1698 VGND.n317 VGND.n306 2.09737
R1699 VGND.n317 VGND.n316 2.09737
R1700 VGND.n426 VGND.n389 2.09737
R1701 VGND.n436 VGND.n389 2.09737
R1702 VGND.n240 VGND.n232 2.09113
R1703 VGND.n481 VGND.n443 2.09113
R1704 VGND.n719 VGND.n681 2.09113
R1705 VGND.n813 VGND.n805 2.09113
R1706 VGND.n992 VGND.n954 2.09113
R1707 VGND.n939 VGND.n901 2.09113
R1708 VGND.n314 VGND.n306 2.09113
R1709 VGND.n426 VGND.n388 2.09113
R1710 VGND.n237 VGND.n236 1.93989
R1711 VGND.n484 VGND.n482 1.93989
R1712 VGND.n722 VGND.n720 1.93989
R1713 VGND.n810 VGND.n809 1.93989
R1714 VGND.n995 VGND.n993 1.93989
R1715 VGND.n942 VGND.n940 1.93989
R1716 VGND.n311 VGND.n310 1.93989
R1717 VGND.n429 VGND.n427 1.93989
R1718 VGND.n241 VGND.n240 1.72862
R1719 VGND.n492 VGND.n443 1.72862
R1720 VGND.n730 VGND.n681 1.72862
R1721 VGND.n814 VGND.n813 1.72862
R1722 VGND.n1003 VGND.n954 1.72862
R1723 VGND.n950 VGND.n901 1.72862
R1724 VGND.n315 VGND.n314 1.72862
R1725 VGND.n437 VGND.n388 1.72862
R1726 VGND.n197 VGND.n196 1.24162
R1727 VGND.n126 VGND.n125 1.24162
R1728 VGND.n654 VGND.n653 1.24162
R1729 VGND.n680 VGND.n679 1.24162
R1730 VGND.n900 VGND.n899 1.24162
R1731 VGND.n874 VGND.n873 1.24162
R1732 VGND.n521 VGND.n520 1.24162
R1733 VGND.n27 VGND.n26 1.24162
R1734 VGND.n738 VGND.t421 1.00615
R1735 VGND.n244 VGND.n231 0.970197
R1736 VGND.n245 VGND.n230 0.970197
R1737 VGND.n239 VGND.n238 0.970197
R1738 VGND.n483 VGND.n446 0.970197
R1739 VGND.n490 VGND.n489 0.970197
R1740 VGND.n480 VGND.n445 0.970197
R1741 VGND.n721 VGND.n684 0.970197
R1742 VGND.n728 VGND.n727 0.970197
R1743 VGND.n718 VGND.n683 0.970197
R1744 VGND.n817 VGND.n804 0.970197
R1745 VGND.n818 VGND.n803 0.970197
R1746 VGND.n812 VGND.n811 0.970197
R1747 VGND.n994 VGND.n957 0.970197
R1748 VGND.n1001 VGND.n1000 0.970197
R1749 VGND.n991 VGND.n956 0.970197
R1750 VGND.n941 VGND.n904 0.970197
R1751 VGND.n948 VGND.n947 0.970197
R1752 VGND.n938 VGND.n903 0.970197
R1753 VGND.n318 VGND.n305 0.970197
R1754 VGND.n319 VGND.n304 0.970197
R1755 VGND.n313 VGND.n312 0.970197
R1756 VGND.n428 VGND.n391 0.970197
R1757 VGND.n435 VGND.n434 0.970197
R1758 VGND.n425 VGND.n390 0.970197
R1759 VGND.n227 VGND.n225 0.927299
R1760 VGND.n476 VGND.n474 0.927299
R1761 VGND.n714 VGND.n712 0.927299
R1762 VGND.n800 VGND.n798 0.927299
R1763 VGND.n987 VGND.n985 0.927299
R1764 VGND.n934 VGND.n932 0.927299
R1765 VGND.n301 VGND.n299 0.927299
R1766 VGND.n421 VGND.n419 0.927299
R1767 VGND.n1092 VGND.n1 0.8465
R1768 VGND.n1093 VGND.n1092 0.8465
R1769 VGND.n253 VGND.n252 0.846456
R1770 VGND.n441 VGND.n83 0.846456
R1771 VGND.n1035 VGND.n1034 0.846456
R1772 VGND.n834 VGND.n833 0.846456
R1773 VGND.n1048 VGND.n1047 0.846456
R1774 VGND.n1076 VGND.n1075 0.846456
R1775 VGND.n327 VGND.n326 0.846456
R1776 VGND.n386 VGND.n385 0.846456
R1777 VGND.n628 VGND.n580 0.721167
R1778 VGND.n213 VGND.n211 0.690273
R1779 VGND.n461 VGND.n459 0.690273
R1780 VGND.n699 VGND.n697 0.690273
R1781 VGND.n786 VGND.n784 0.690273
R1782 VGND.n972 VGND.n970 0.690273
R1783 VGND.n919 VGND.n917 0.690273
R1784 VGND.n287 VGND.n285 0.690273
R1785 VGND.n406 VGND.n404 0.690273
R1786 VGND.n225 VGND.n214 0.60675
R1787 VGND.n474 VGND.n463 0.60675
R1788 VGND.n712 VGND.n701 0.60675
R1789 VGND.n798 VGND.n787 0.60675
R1790 VGND.n985 VGND.n974 0.60675
R1791 VGND.n932 VGND.n921 0.60675
R1792 VGND.n299 VGND.n288 0.60675
R1793 VGND.n419 VGND.n408 0.60675
R1794 VGND.n1063 VGND.n59 0.5455
R1795 VGND.n733 VGND.n627 0.5455
R1796 VGND.n1016 VGND.n1006 0.5455
R1797 VGND.n953 VGND.n848 0.5455
R1798 VGND.n771 VGND.n770 0.5455
R1799 VGND.n523 VGND.n522 0.5455
R1800 VGND.n358 VGND.n0 0.5455
R1801 VGND.n1091 VGND.n1090 0.5455
R1802 VGND.n225 VGND.n219 0.516045
R1803 VGND.n474 VGND.n468 0.516045
R1804 VGND.n712 VGND.n706 0.516045
R1805 VGND.n798 VGND.n792 0.516045
R1806 VGND.n985 VGND.n979 0.516045
R1807 VGND.n932 VGND.n926 0.516045
R1808 VGND.n299 VGND.n293 0.516045
R1809 VGND.n419 VGND.n413 0.516045
R1810 VGND.n215 VGND.n214 0.454213
R1811 VGND.n464 VGND.n463 0.454213
R1812 VGND.n702 VGND.n701 0.454213
R1813 VGND.n788 VGND.n787 0.454213
R1814 VGND.n975 VGND.n974 0.454213
R1815 VGND.n922 VGND.n921 0.454213
R1816 VGND.n289 VGND.n288 0.454213
R1817 VGND.n409 VGND.n408 0.454213
R1818 VGND.n258 VGND.n168 0.376971
R1819 VGND.n537 VGND.n85 0.376971
R1820 VGND.n560 VGND.n554 0.376971
R1821 VGND.n828 VGND.n602 0.376971
R1822 VGND.n45 VGND.n39 0.376971
R1823 VGND.n332 VGND.n142 0.376971
R1824 VGND.n376 VGND.n375 0.376971
R1825 VGND.n242 VGND.n241 0.363
R1826 VGND.n492 VGND.n491 0.363
R1827 VGND.n730 VGND.n729 0.363
R1828 VGND.n815 VGND.n814 0.363
R1829 VGND.n1003 VGND.n1002 0.363
R1830 VGND.n950 VGND.n949 0.363
R1831 VGND.n316 VGND.n315 0.363
R1832 VGND.n437 VGND.n436 0.363
R1833 VGND.n222 VGND.n214 0.347226
R1834 VGND.n471 VGND.n463 0.347226
R1835 VGND.n709 VGND.n701 0.347226
R1836 VGND.n795 VGND.n787 0.347226
R1837 VGND.n982 VGND.n974 0.347226
R1838 VGND.n929 VGND.n921 0.347226
R1839 VGND.n296 VGND.n288 0.347226
R1840 VGND.n416 VGND.n408 0.347226
R1841 VGND.n240 VGND.n239 0.344944
R1842 VGND.n244 VGND.n243 0.344944
R1843 VGND.n445 VGND.n443 0.344944
R1844 VGND.n446 VGND.n444 0.344944
R1845 VGND.n683 VGND.n681 0.344944
R1846 VGND.n684 VGND.n682 0.344944
R1847 VGND.n813 VGND.n812 0.344944
R1848 VGND.n817 VGND.n816 0.344944
R1849 VGND.n956 VGND.n954 0.344944
R1850 VGND.n957 VGND.n955 0.344944
R1851 VGND.n903 VGND.n901 0.344944
R1852 VGND.n904 VGND.n902 0.344944
R1853 VGND.n314 VGND.n313 0.344944
R1854 VGND.n318 VGND.n317 0.344944
R1855 VGND.n390 VGND.n388 0.344944
R1856 VGND.n391 VGND.n389 0.344944
R1857 VGND.n216 VGND.n215 0.319807
R1858 VGND.n465 VGND.n464 0.319807
R1859 VGND.n703 VGND.n702 0.319807
R1860 VGND.n789 VGND.n788 0.319807
R1861 VGND.n976 VGND.n975 0.319807
R1862 VGND.n923 VGND.n922 0.319807
R1863 VGND.n290 VGND.n289 0.319807
R1864 VGND.n410 VGND.n409 0.319807
R1865 VGND.n219 VGND.n218 0.291342
R1866 VGND.n468 VGND.n467 0.291342
R1867 VGND.n706 VGND.n705 0.291342
R1868 VGND.n792 VGND.n791 0.291342
R1869 VGND.n979 VGND.n978 0.291342
R1870 VGND.n926 VGND.n925 0.291342
R1871 VGND.n293 VGND.n292 0.291342
R1872 VGND.n413 VGND.n412 0.291342
R1873 VGND.n222 VGND.n219 0.22669
R1874 VGND.n471 VGND.n468 0.22669
R1875 VGND.n709 VGND.n706 0.22669
R1876 VGND.n795 VGND.n792 0.22669
R1877 VGND.n982 VGND.n979 0.22669
R1878 VGND.n929 VGND.n926 0.22669
R1879 VGND.n296 VGND.n293 0.22669
R1880 VGND.n416 VGND.n413 0.22669
R1881 VGND.n250 VGND.n213 0.216409
R1882 VGND.n462 VGND.n461 0.216409
R1883 VGND.n700 VGND.n699 0.216409
R1884 VGND.n823 VGND.n786 0.216409
R1885 VGND.n973 VGND.n972 0.216409
R1886 VGND.n920 VGND.n919 0.216409
R1887 VGND.n324 VGND.n287 0.216409
R1888 VGND.n407 VGND.n406 0.216409
R1889 VGND.n249 VGND.n227 0.210727
R1890 VGND.n477 VGND.n476 0.210727
R1891 VGND.n715 VGND.n714 0.210727
R1892 VGND.n822 VGND.n800 0.210727
R1893 VGND.n988 VGND.n987 0.210727
R1894 VGND.n935 VGND.n934 0.210727
R1895 VGND.n323 VGND.n301 0.210727
R1896 VGND.n422 VGND.n421 0.210727
R1897 VGND VGND.n1095 0.198859
R1898 VGND.n252 VGND.n251 0.158833
R1899 VGND.n442 VGND.n441 0.158833
R1900 VGND.n1035 VGND.n556 0.158833
R1901 VGND.n834 VGND.n824 0.158833
R1902 VGND.n1048 VGND.n74 0.158833
R1903 VGND.n1076 VGND.n41 0.158833
R1904 VGND.n326 VGND.n325 0.158833
R1905 VGND.n387 VGND.n386 0.158833
R1906 VGND.n220 VGND.n219 0.158238
R1907 VGND.n469 VGND.n468 0.158238
R1908 VGND.n707 VGND.n706 0.158238
R1909 VGND.n793 VGND.n792 0.158238
R1910 VGND.n980 VGND.n979 0.158238
R1911 VGND.n927 VGND.n926 0.158238
R1912 VGND.n294 VGND.n293 0.158238
R1913 VGND.n414 VGND.n413 0.158238
R1914 VGND.n522 VGND 0.149613
R1915 VGND VGND.n1091 0.14291
R1916 VGND.n521 VGND.n495 0.142507
R1917 VGND.n272 VGND.n27 0.142507
R1918 VGND.n198 VGND.n197 0.142507
R1919 VGND.n440 VGND.n126 0.1417
R1920 VGND.n237 VGND.n232 0.135283
R1921 VGND.n242 VGND.n230 0.135283
R1922 VGND.n482 VGND.n481 0.135283
R1923 VGND.n491 VGND.n490 0.135283
R1924 VGND.n720 VGND.n719 0.135283
R1925 VGND.n729 VGND.n728 0.135283
R1926 VGND.n810 VGND.n805 0.135283
R1927 VGND.n815 VGND.n803 0.135283
R1928 VGND.n993 VGND.n992 0.135283
R1929 VGND.n1002 VGND.n1001 0.135283
R1930 VGND.n940 VGND.n939 0.135283
R1931 VGND.n949 VGND.n948 0.135283
R1932 VGND.n311 VGND.n306 0.135283
R1933 VGND.n316 VGND.n304 0.135283
R1934 VGND.n427 VGND.n426 0.135283
R1935 VGND.n436 VGND.n435 0.135283
R1936 VGND VGND.n59 0.133711
R1937 VGND.n177 VGND.n176 0.120292
R1938 VGND.n177 VGND.n172 0.120292
R1939 VGND.n195 VGND.n173 0.120292
R1940 VGND.n190 VGND.n173 0.120292
R1941 VGND.n190 VGND.n189 0.120292
R1942 VGND.n189 VGND.n184 0.120292
R1943 VGND.n185 VGND.n184 0.120292
R1944 VGND.n106 VGND.n105 0.120292
R1945 VGND.n106 VGND.n101 0.120292
R1946 VGND.n124 VGND.n102 0.120292
R1947 VGND.n119 VGND.n102 0.120292
R1948 VGND.n119 VGND.n118 0.120292
R1949 VGND.n118 VGND.n113 0.120292
R1950 VGND.n114 VGND.n113 0.120292
R1951 VGND.n634 VGND.n633 0.120292
R1952 VGND.n634 VGND.n629 0.120292
R1953 VGND.n652 VGND.n630 0.120292
R1954 VGND.n647 VGND.n630 0.120292
R1955 VGND.n647 VGND.n646 0.120292
R1956 VGND.n646 VGND.n641 0.120292
R1957 VGND.n642 VGND.n641 0.120292
R1958 VGND.n660 VGND.n659 0.120292
R1959 VGND.n660 VGND.n655 0.120292
R1960 VGND.n678 VGND.n656 0.120292
R1961 VGND.n673 VGND.n656 0.120292
R1962 VGND.n673 VGND.n672 0.120292
R1963 VGND.n672 VGND.n667 0.120292
R1964 VGND.n668 VGND.n667 0.120292
R1965 VGND.n880 VGND.n879 0.120292
R1966 VGND.n880 VGND.n875 0.120292
R1967 VGND.n898 VGND.n876 0.120292
R1968 VGND.n893 VGND.n876 0.120292
R1969 VGND.n893 VGND.n892 0.120292
R1970 VGND.n892 VGND.n887 0.120292
R1971 VGND.n888 VGND.n887 0.120292
R1972 VGND.n854 VGND.n853 0.120292
R1973 VGND.n854 VGND.n849 0.120292
R1974 VGND.n872 VGND.n850 0.120292
R1975 VGND.n867 VGND.n850 0.120292
R1976 VGND.n867 VGND.n866 0.120292
R1977 VGND.n866 VGND.n861 0.120292
R1978 VGND.n862 VGND.n861 0.120292
R1979 VGND.n501 VGND.n500 0.120292
R1980 VGND.n501 VGND.n496 0.120292
R1981 VGND.n519 VGND.n497 0.120292
R1982 VGND.n514 VGND.n497 0.120292
R1983 VGND.n514 VGND.n513 0.120292
R1984 VGND.n513 VGND.n508 0.120292
R1985 VGND.n509 VGND.n508 0.120292
R1986 VGND.n7 VGND.n6 0.120292
R1987 VGND.n7 VGND.n2 0.120292
R1988 VGND.n25 VGND.n3 0.120292
R1989 VGND.n20 VGND.n3 0.120292
R1990 VGND.n20 VGND.n19 0.120292
R1991 VGND.n19 VGND.n14 0.120292
R1992 VGND.n15 VGND.n14 0.120292
R1993 VGND.n196 VGND.n172 0.112479
R1994 VGND.n125 VGND.n101 0.112479
R1995 VGND.n653 VGND.n629 0.112479
R1996 VGND.n679 VGND.n655 0.112479
R1997 VGND.n899 VGND.n875 0.112479
R1998 VGND.n873 VGND.n849 0.112479
R1999 VGND.n520 VGND.n496 0.112479
R2000 VGND.n26 VGND.n2 0.112479
R2001 VGND.n251 VGND.n250 0.09425
R2002 VGND.n462 VGND.n442 0.09425
R2003 VGND.n700 VGND.n556 0.09425
R2004 VGND.n824 VGND.n823 0.09425
R2005 VGND.n973 VGND.n74 0.09425
R2006 VGND.n920 VGND.n41 0.09425
R2007 VGND.n325 VGND.n324 0.09425
R2008 VGND.n407 VGND.n387 0.09425
R2009 VGND.n495 VGND 0.0941643
R2010 VGND.n272 VGND 0.0941643
R2011 VGND.n198 VGND 0.0941643
R2012 VGND VGND.n440 0.0936321
R2013 VGND.n218 VGND.n217 0.0714406
R2014 VGND.n467 VGND.n466 0.0714406
R2015 VGND.n705 VGND.n704 0.0714406
R2016 VGND.n791 VGND.n790 0.0714406
R2017 VGND.n978 VGND.n977 0.0714406
R2018 VGND.n925 VGND.n924 0.0714406
R2019 VGND.n292 VGND.n291 0.0714406
R2020 VGND.n412 VGND.n411 0.0714406
R2021 VGND.n628 VGND 0.0610165
R2022 VGND.n176 VGND 0.0603958
R2023 VGND.n105 VGND 0.0603958
R2024 VGND.n633 VGND 0.0603958
R2025 VGND.n659 VGND 0.0603958
R2026 VGND.n879 VGND 0.0603958
R2027 VGND.n853 VGND 0.0603958
R2028 VGND.n500 VGND 0.0603958
R2029 VGND.n6 VGND 0.0603958
R2030 VGND.n200 VGND.n199 0.0584812
R2031 VGND.n494 VGND.n493 0.0584812
R2032 VGND.n732 VGND.n731 0.0584812
R2033 VGND.n773 VGND.n772 0.0584812
R2034 VGND.n1005 VGND.n1004 0.0584812
R2035 VGND.n952 VGND.n951 0.0584812
R2036 VGND.n274 VGND.n273 0.0584812
R2037 VGND.n439 VGND.n438 0.0584812
R2038 VGND.n522 VGND.n521 0.0582429
R2039 VGND.n1091 VGND.n27 0.0582429
R2040 VGND.n197 VGND.n59 0.0582429
R2041 VGND.n126 VGND.n0 0.0579148
R2042 VGND.n199 VGND 0.0520484
R2043 VGND.n494 VGND 0.0520484
R2044 VGND.n732 VGND 0.0520484
R2045 VGND.n772 VGND 0.0520484
R2046 VGND.n1005 VGND 0.0520484
R2047 VGND.n952 VGND 0.0520484
R2048 VGND.n273 VGND 0.0520484
R2049 VGND.n439 VGND 0.0520484
R2050 VGND.n1 VGND 0.0503372
R2051 VGND VGND.n359 0.0459545
R2052 VGND VGND.n1064 0.0459545
R2053 VGND.n1062 VGND 0.0459545
R2054 VGND.n769 VGND 0.0459545
R2055 VGND.n618 VGND 0.0459545
R2056 VGND.n626 VGND 0.0459545
R2057 VGND VGND.n1017 0.0459545
R2058 VGND.n1015 VGND 0.0459545
R2059 VGND VGND.n581 0.0459545
R2060 VGND.n847 VGND 0.0459545
R2061 VGND VGND.n734 0.0459545
R2062 VGND VGND.n28 0.0459545
R2063 VGND VGND.n100 0.0459545
R2064 VGND VGND.n524 0.0459545
R2065 VGND.n357 VGND 0.0459545
R2066 VGND.n1089 VGND 0.0459545
R2067 VGND.n241 VGND.n200 0.0455
R2068 VGND.n493 VGND.n492 0.0455
R2069 VGND.n731 VGND.n730 0.0455
R2070 VGND.n814 VGND.n773 0.0455
R2071 VGND.n1004 VGND.n1003 0.0455
R2072 VGND.n951 VGND.n950 0.0455
R2073 VGND.n315 VGND.n274 0.0455
R2074 VGND.n438 VGND.n437 0.0455
R2075 VGND.n206 VGND.n202 0.0429342
R2076 VGND.n207 VGND.n206 0.0429342
R2077 VGND.n208 VGND.n207 0.0429342
R2078 VGND.n208 VGND.n201 0.0429342
R2079 VGND.n454 VGND.n450 0.0429342
R2080 VGND.n455 VGND.n454 0.0429342
R2081 VGND.n456 VGND.n455 0.0429342
R2082 VGND.n456 VGND.n449 0.0429342
R2083 VGND.n692 VGND.n688 0.0429342
R2084 VGND.n693 VGND.n692 0.0429342
R2085 VGND.n694 VGND.n693 0.0429342
R2086 VGND.n694 VGND.n687 0.0429342
R2087 VGND.n779 VGND.n775 0.0429342
R2088 VGND.n780 VGND.n779 0.0429342
R2089 VGND.n781 VGND.n780 0.0429342
R2090 VGND.n781 VGND.n774 0.0429342
R2091 VGND.n965 VGND.n961 0.0429342
R2092 VGND.n966 VGND.n965 0.0429342
R2093 VGND.n967 VGND.n966 0.0429342
R2094 VGND.n967 VGND.n960 0.0429342
R2095 VGND.n912 VGND.n908 0.0429342
R2096 VGND.n913 VGND.n912 0.0429342
R2097 VGND.n914 VGND.n913 0.0429342
R2098 VGND.n914 VGND.n907 0.0429342
R2099 VGND.n280 VGND.n276 0.0429342
R2100 VGND.n281 VGND.n280 0.0429342
R2101 VGND.n282 VGND.n281 0.0429342
R2102 VGND.n282 VGND.n275 0.0429342
R2103 VGND.n399 VGND.n395 0.0429342
R2104 VGND.n400 VGND.n399 0.0429342
R2105 VGND.n401 VGND.n400 0.0429342
R2106 VGND.n401 VGND.n394 0.0429342
R2107 VGND.n204 VGND.n203 0.0389615
R2108 VGND.n452 VGND.n451 0.0389615
R2109 VGND.n690 VGND.n689 0.0389615
R2110 VGND.n777 VGND.n776 0.0389615
R2111 VGND.n963 VGND.n962 0.0389615
R2112 VGND.n910 VGND.n909 0.0389615
R2113 VGND.n278 VGND.n277 0.0389615
R2114 VGND.n397 VGND.n396 0.0389615
R2115 VGND.n211 VGND.n201 0.0340526
R2116 VGND.n459 VGND.n449 0.0340526
R2117 VGND.n697 VGND.n687 0.0340526
R2118 VGND.n784 VGND.n774 0.0340526
R2119 VGND.n970 VGND.n960 0.0340526
R2120 VGND.n917 VGND.n907 0.0340526
R2121 VGND.n285 VGND.n275 0.0340526
R2122 VGND.n404 VGND.n394 0.0340526
R2123 VGND.n359 VGND 0.0338333
R2124 VGND.n1064 VGND 0.0338333
R2125 VGND.n1062 VGND 0.0338333
R2126 VGND.n769 VGND 0.0338333
R2127 VGND.n618 VGND 0.0338333
R2128 VGND.n626 VGND 0.0338333
R2129 VGND.n1017 VGND 0.0338333
R2130 VGND.n1015 VGND 0.0338333
R2131 VGND.n581 VGND 0.0338333
R2132 VGND.n847 VGND 0.0338333
R2133 VGND.n734 VGND 0.0338333
R2134 VGND.n28 VGND 0.0338333
R2135 VGND.n100 VGND 0.0338333
R2136 VGND.n524 VGND 0.0338333
R2137 VGND.n357 VGND 0.0338333
R2138 VGND.n1089 VGND 0.0338333
R2139 VGND.n219 VGND.n216 0.0289653
R2140 VGND.n468 VGND.n465 0.0289653
R2141 VGND.n706 VGND.n703 0.0289653
R2142 VGND.n792 VGND.n789 0.0289653
R2143 VGND.n979 VGND.n976 0.0289653
R2144 VGND.n926 VGND.n923 0.0289653
R2145 VGND.n293 VGND.n290 0.0289653
R2146 VGND.n413 VGND.n410 0.0289653
R2147 VGND.n1094 VGND.n0 0.0265369
R2148 VGND.n185 VGND 0.0226354
R2149 VGND.n114 VGND 0.0226354
R2150 VGND.n642 VGND 0.0226354
R2151 VGND.n668 VGND 0.0226354
R2152 VGND.n888 VGND 0.0226354
R2153 VGND.n862 VGND 0.0226354
R2154 VGND.n509 VGND 0.0226354
R2155 VGND.n15 VGND 0.0226354
R2156 VGND.n1094 VGND.n1093 0.0101424
R2157 VGND.n1095 VGND.n1094 0.0101424
R2158 VGND.n196 VGND.n195 0.0083125
R2159 VGND.n125 VGND.n124 0.0083125
R2160 VGND.n653 VGND.n652 0.0083125
R2161 VGND.n679 VGND.n678 0.0083125
R2162 VGND.n899 VGND.n898 0.0083125
R2163 VGND.n873 VGND.n872 0.0083125
R2164 VGND.n520 VGND.n519 0.0083125
R2165 VGND.n26 VGND.n25 0.0083125
R2166 VGND.n204 VGND.n202 0.00773684
R2167 VGND.n452 VGND.n450 0.00773684
R2168 VGND.n690 VGND.n688 0.00773684
R2169 VGND.n777 VGND.n775 0.00773684
R2170 VGND.n963 VGND.n961 0.00773684
R2171 VGND.n910 VGND.n908 0.00773684
R2172 VGND.n278 VGND.n276 0.00773684
R2173 VGND.n397 VGND.n395 0.00773684
R2174 VGND.n250 VGND.n249 0.00618182
R2175 VGND.n477 VGND.n462 0.00618182
R2176 VGND.n715 VGND.n700 0.00618182
R2177 VGND.n823 VGND.n822 0.00618182
R2178 VGND.n988 VGND.n973 0.00618182
R2179 VGND.n935 VGND.n920 0.00618182
R2180 VGND.n324 VGND.n323 0.00618182
R2181 VGND.n422 VGND.n407 0.00618182
R2182 VGND.n1092 VGND 0.00553571
R2183 VGND.n953 VGND.n952 0.00544203
R2184 VGND.n1006 VGND.n1005 0.00544203
R2185 VGND.n772 VGND.n771 0.00544203
R2186 VGND.n733 VGND.n732 0.00544203
R2187 VGND.n495 VGND.n494 0.00544203
R2188 VGND.n440 VGND.n439 0.00544203
R2189 VGND.n273 VGND.n272 0.00544203
R2190 VGND.n199 VGND.n198 0.00544203
R2191 VGND.n1006 VGND.n580 0.00167117
R2192 VGND.n251 VGND.n200 0.00154167
R2193 VGND.n493 VGND.n442 0.00154167
R2194 VGND.n731 VGND.n556 0.00154167
R2195 VGND.n824 VGND.n773 0.00154167
R2196 VGND.n1004 VGND.n74 0.00154167
R2197 VGND.n951 VGND.n41 0.00154167
R2198 VGND.n325 VGND.n274 0.00154167
R2199 VGND.n438 VGND.n387 0.00154167
R2200 VGND VGND.n1 0.000955654
R2201 VGND VGND.n628 0.000891578
R2202 VGND.n953 VGND.n900 0.0008453
R2203 VGND.n771 VGND.n733 0.000777664
R2204 VGND.n680 VGND 0.000749186
R2205 VGND.n654 VGND 0.000749186
R2206 VGND.n733 VGND.n680 0.000702908
R2207 VGND.n1006 VGND.n953 0.000635272
R2208 VGND.n900 VGND.n874 0.000635272
R2209 VGND.n874 VGND 0.000613914
R2210 VGND VGND.n654 0.000528478
R2211 VPWR.n174 VPWR.n173 18810
R2212 VPWR.n253 VPWR.n252 18810
R2213 VPWR.n93 VPWR.n92 18810
R2214 VPWR.n14 VPWR.n13 18810
R2215 VPWR.n455 VPWR.n454 18810
R2216 VPWR.n374 VPWR.n373 18810
R2217 VPWR.n617 VPWR.n616 18810
R2218 VPWR.n536 VPWR.n535 18810
R2219 VPWR.n175 VPWR.n174 18786.2
R2220 VPWR.n175 VPWR.n166 18786.2
R2221 VPWR.n254 VPWR.n253 18786.2
R2222 VPWR.n254 VPWR.n245 18786.2
R2223 VPWR.n94 VPWR.n93 18786.2
R2224 VPWR.n94 VPWR.n85 18786.2
R2225 VPWR.n15 VPWR.n14 18786.2
R2226 VPWR.n15 VPWR.n6 18786.2
R2227 VPWR.n456 VPWR.n455 18786.2
R2228 VPWR.n456 VPWR.n447 18786.2
R2229 VPWR.n375 VPWR.n374 18786.2
R2230 VPWR.n375 VPWR.n366 18786.2
R2231 VPWR.n618 VPWR.n617 18786.2
R2232 VPWR.n618 VPWR.n609 18786.2
R2233 VPWR.n537 VPWR.n536 18786.2
R2234 VPWR.n537 VPWR.n528 18786.2
R2235 VPWR.n173 VPWR.n166 18667.5
R2236 VPWR.n252 VPWR.n245 18667.5
R2237 VPWR.n92 VPWR.n85 18667.5
R2238 VPWR.n13 VPWR.n6 18667.5
R2239 VPWR.n454 VPWR.n447 18667.5
R2240 VPWR.n373 VPWR.n366 18667.5
R2241 VPWR.n616 VPWR.n609 18667.5
R2242 VPWR.n535 VPWR.n528 18667.5
R2243 VPWR.n176 VPWR.n164 7334.54
R2244 VPWR.n255 VPWR.n243 7334.54
R2245 VPWR.n95 VPWR.n83 7334.54
R2246 VPWR.n16 VPWR.n4 7334.54
R2247 VPWR.n457 VPWR.n445 7334.54
R2248 VPWR.n376 VPWR.n364 7334.54
R2249 VPWR.n619 VPWR.n607 7334.54
R2250 VPWR.n538 VPWR.n526 7334.54
R2251 VPWR.n172 VPWR.n165 7332.73
R2252 VPWR.n251 VPWR.n244 7332.73
R2253 VPWR.n91 VPWR.n84 7332.73
R2254 VPWR.n12 VPWR.n5 7332.73
R2255 VPWR.n453 VPWR.n446 7332.73
R2256 VPWR.n372 VPWR.n365 7332.73
R2257 VPWR.n615 VPWR.n608 7332.73
R2258 VPWR.n534 VPWR.n527 7332.73
R2259 VPWR.n176 VPWR.n165 7312.73
R2260 VPWR.n255 VPWR.n244 7312.73
R2261 VPWR.n95 VPWR.n84 7312.73
R2262 VPWR.n16 VPWR.n5 7312.73
R2263 VPWR.n457 VPWR.n446 7312.73
R2264 VPWR.n376 VPWR.n365 7312.73
R2265 VPWR.n619 VPWR.n608 7312.73
R2266 VPWR.n538 VPWR.n527 7312.73
R2267 VPWR.n172 VPWR.n164 7300
R2268 VPWR.n251 VPWR.n243 7300
R2269 VPWR.n91 VPWR.n83 7300
R2270 VPWR.n12 VPWR.n4 7300
R2271 VPWR.n453 VPWR.n445 7300
R2272 VPWR.n372 VPWR.n364 7300
R2273 VPWR.n615 VPWR.n607 7300
R2274 VPWR.n534 VPWR.n526 7300
R2275 VPWR.n227 VPWR.n225 4136.47
R2276 VPWR.n234 VPWR.n232 4136.47
R2277 VPWR.n306 VPWR.n304 4136.47
R2278 VPWR.n313 VPWR.n311 4136.47
R2279 VPWR.n67 VPWR.n65 4136.47
R2280 VPWR.n74 VPWR.n72 4136.47
R2281 VPWR.n146 VPWR.n144 4136.47
R2282 VPWR.n153 VPWR.n151 4136.47
R2283 VPWR.n403 VPWR.n401 4136.47
R2284 VPWR.n410 VPWR.n408 4136.47
R2285 VPWR.n323 VPWR.n321 4136.47
R2286 VPWR.n330 VPWR.n328 4136.47
R2287 VPWR.n565 VPWR.n563 4136.47
R2288 VPWR.n572 VPWR.n570 4136.47
R2289 VPWR.n485 VPWR.n483 4136.47
R2290 VPWR.n492 VPWR.n490 4136.47
R2291 VPWR.n227 VPWR.n224 2068.24
R2292 VPWR.n234 VPWR.n231 2068.24
R2293 VPWR.n306 VPWR.n303 2068.24
R2294 VPWR.n313 VPWR.n310 2068.24
R2295 VPWR.n67 VPWR.n64 2068.24
R2296 VPWR.n74 VPWR.n71 2068.24
R2297 VPWR.n146 VPWR.n143 2068.24
R2298 VPWR.n153 VPWR.n150 2068.24
R2299 VPWR.n403 VPWR.n400 2068.24
R2300 VPWR.n410 VPWR.n407 2068.24
R2301 VPWR.n323 VPWR.n320 2068.24
R2302 VPWR.n330 VPWR.n327 2068.24
R2303 VPWR.n565 VPWR.n562 2068.24
R2304 VPWR.n572 VPWR.n569 2068.24
R2305 VPWR.n485 VPWR.n482 2068.24
R2306 VPWR.n492 VPWR.n489 2068.24
R2307 VPWR.n170 VPWR.n168 781.188
R2308 VPWR.n249 VPWR.n247 781.188
R2309 VPWR.n89 VPWR.n87 781.188
R2310 VPWR.n10 VPWR.n8 781.188
R2311 VPWR.n451 VPWR.n449 781.188
R2312 VPWR.n370 VPWR.n368 781.188
R2313 VPWR.n613 VPWR.n611 781.188
R2314 VPWR.n532 VPWR.n530 781.188
R2315 VPWR.n178 VPWR.n162 779.442
R2316 VPWR.n257 VPWR.n241 779.442
R2317 VPWR.n97 VPWR.n81 779.442
R2318 VPWR.n18 VPWR.n2 779.442
R2319 VPWR.n459 VPWR.n443 779.442
R2320 VPWR.n378 VPWR.n362 779.442
R2321 VPWR.n621 VPWR.n605 779.442
R2322 VPWR.n540 VPWR.n524 779.442
R2323 VPWR.n177 VPWR.n163 779.056
R2324 VPWR.n256 VPWR.n242 779.056
R2325 VPWR.n96 VPWR.n82 779.056
R2326 VPWR.n17 VPWR.n3 779.056
R2327 VPWR.n458 VPWR.n444 779.056
R2328 VPWR.n377 VPWR.n363 779.056
R2329 VPWR.n620 VPWR.n606 779.056
R2330 VPWR.n539 VPWR.n525 779.056
R2331 VPWR.n171 VPWR.n167 778.668
R2332 VPWR.n250 VPWR.n246 778.668
R2333 VPWR.n90 VPWR.n86 778.668
R2334 VPWR.n11 VPWR.n7 778.668
R2335 VPWR.n452 VPWR.n448 778.668
R2336 VPWR.n371 VPWR.n367 778.668
R2337 VPWR.n614 VPWR.n610 778.668
R2338 VPWR.n533 VPWR.n529 778.668
R2339 VPWR.t143 VPWR.t242 478.712
R2340 VPWR.t149 VPWR.t143 478.712
R2341 VPWR.t153 VPWR.t149 478.712
R2342 VPWR.t141 VPWR.t153 478.712
R2343 VPWR.t139 VPWR.t141 478.712
R2344 VPWR.t145 VPWR.t147 478.712
R2345 VPWR.t147 VPWR.t151 478.712
R2346 VPWR.t151 VPWR.t137 478.712
R2347 VPWR.t137 VPWR.t155 478.712
R2348 VPWR.t155 VPWR.t239 478.712
R2349 VPWR.t164 VPWR.t230 478.712
R2350 VPWR.t168 VPWR.t164 478.712
R2351 VPWR.t174 VPWR.t168 478.712
R2352 VPWR.t160 VPWR.t174 478.712
R2353 VPWR.t178 VPWR.t160 478.712
R2354 VPWR.t162 VPWR.t166 478.712
R2355 VPWR.t166 VPWR.t172 478.712
R2356 VPWR.t172 VPWR.t170 478.712
R2357 VPWR.t170 VPWR.t176 478.712
R2358 VPWR.t176 VPWR.t236 478.712
R2359 VPWR.t92 VPWR.t248 478.712
R2360 VPWR.t94 VPWR.t92 478.712
R2361 VPWR.t102 VPWR.t94 478.712
R2362 VPWR.t100 VPWR.t102 478.712
R2363 VPWR.t106 VPWR.t100 478.712
R2364 VPWR.t108 VPWR.t90 478.712
R2365 VPWR.t90 VPWR.t98 478.712
R2366 VPWR.t98 VPWR.t96 478.712
R2367 VPWR.t96 VPWR.t104 478.712
R2368 VPWR.t104 VPWR.t257 478.712
R2369 VPWR.t209 VPWR.t260 478.712
R2370 VPWR.t193 VPWR.t209 478.712
R2371 VPWR.t197 VPWR.t193 478.712
R2372 VPWR.t201 VPWR.t197 478.712
R2373 VPWR.t207 VPWR.t201 478.712
R2374 VPWR.t205 VPWR.t211 478.712
R2375 VPWR.t211 VPWR.t195 478.712
R2376 VPWR.t195 VPWR.t199 478.712
R2377 VPWR.t199 VPWR.t203 478.712
R2378 VPWR.t203 VPWR.t251 478.712
R2379 VPWR.t65 VPWR.t224 478.712
R2380 VPWR.t69 VPWR.t65 478.712
R2381 VPWR.t73 VPWR.t69 478.712
R2382 VPWR.t61 VPWR.t73 478.712
R2383 VPWR.t59 VPWR.t61 478.712
R2384 VPWR.t67 VPWR.t63 478.712
R2385 VPWR.t63 VPWR.t71 478.712
R2386 VPWR.t71 VPWR.t57 478.712
R2387 VPWR.t57 VPWR.t55 478.712
R2388 VPWR.t55 VPWR.t245 478.712
R2389 VPWR.t285 VPWR.t227 478.712
R2390 VPWR.t283 VPWR.t285 478.712
R2391 VPWR.t289 VPWR.t283 478.712
R2392 VPWR.t277 VPWR.t289 478.712
R2393 VPWR.t295 VPWR.t277 478.712
R2394 VPWR.t281 VPWR.t279 478.712
R2395 VPWR.t279 VPWR.t287 478.712
R2396 VPWR.t287 VPWR.t291 478.712
R2397 VPWR.t291 VPWR.t293 478.712
R2398 VPWR.t293 VPWR.t233 478.712
R2399 VPWR.t46 VPWR.t269 478.712
R2400 VPWR.t36 VPWR.t46 478.712
R2401 VPWR.t34 VPWR.t36 478.712
R2402 VPWR.t40 VPWR.t34 478.712
R2403 VPWR.t44 VPWR.t40 478.712
R2404 VPWR.t48 VPWR.t32 478.712
R2405 VPWR.t32 VPWR.t30 478.712
R2406 VPWR.t30 VPWR.t38 478.712
R2407 VPWR.t38 VPWR.t42 478.712
R2408 VPWR.t42 VPWR.t266 478.712
R2409 VPWR.t126 VPWR.t263 478.712
R2410 VPWR.t112 VPWR.t126 478.712
R2411 VPWR.t114 VPWR.t112 478.712
R2412 VPWR.t118 VPWR.t114 478.712
R2413 VPWR.t124 VPWR.t118 478.712
R2414 VPWR.t122 VPWR.t110 478.712
R2415 VPWR.t110 VPWR.t128 478.712
R2416 VPWR.t128 VPWR.t116 478.712
R2417 VPWR.t116 VPWR.t120 478.712
R2418 VPWR.t120 VPWR.t254 478.712
R2419 VPWR.n227 VPWR.t190 452.676
R2420 VPWR.t189 VPWR.n225 452.676
R2421 VPWR.n234 VPWR.t29 452.676
R2422 VPWR.t28 VPWR.n232 452.676
R2423 VPWR.n306 VPWR.t133 452.676
R2424 VPWR.t6 VPWR.n304 452.676
R2425 VPWR.n313 VPWR.t309 452.676
R2426 VPWR.t308 VPWR.n311 452.676
R2427 VPWR.n67 VPWR.t184 452.676
R2428 VPWR.t25 VPWR.n65 452.676
R2429 VPWR.n74 VPWR.t132 452.676
R2430 VPWR.t131 VPWR.n72 452.676
R2431 VPWR.n146 VPWR.t86 452.676
R2432 VPWR.t88 VPWR.n144 452.676
R2433 VPWR.n153 VPWR.t180 452.676
R2434 VPWR.t181 VPWR.n151 452.676
R2435 VPWR.n403 VPWR.t213 452.676
R2436 VPWR.t221 VPWR.n401 452.676
R2437 VPWR.n410 VPWR.t310 452.676
R2438 VPWR.t311 VPWR.n408 452.676
R2439 VPWR.n323 VPWR.t76 452.676
R2440 VPWR.t77 VPWR.n321 452.676
R2441 VPWR.n330 VPWR.t273 452.676
R2442 VPWR.t272 VPWR.n328 452.676
R2443 VPWR.n565 VPWR.t22 452.676
R2444 VPWR.t4 VPWR.n563 452.676
R2445 VPWR.n572 VPWR.t9 452.676
R2446 VPWR.t8 VPWR.n570 452.676
R2447 VPWR.n485 VPWR.t134 452.676
R2448 VPWR.t17 VPWR.n483 452.676
R2449 VPWR.n492 VPWR.t158 452.676
R2450 VPWR.t157 VPWR.n490 452.676
R2451 VPWR.n213 VPWR.t1 342.377
R2452 VPWR.n292 VPWR.t130 342.377
R2453 VPWR.n132 VPWR.t307 342.377
R2454 VPWR.n53 VPWR.t192 342.377
R2455 VPWR.n430 VPWR.t215 342.377
R2456 VPWR.n349 VPWR.t15 342.377
R2457 VPWR.n592 VPWR.t183 342.377
R2458 VPWR.n511 VPWR.t24 342.377
R2459 VPWR.n203 VPWR.t27 338.892
R2460 VPWR.n282 VPWR.t301 338.892
R2461 VPWR.n122 VPWR.t306 338.892
R2462 VPWR.n43 VPWR.t82 338.892
R2463 VPWR.n420 VPWR.t218 338.892
R2464 VPWR.n339 VPWR.t51 338.892
R2465 VPWR.n582 VPWR.t185 338.892
R2466 VPWR.n501 VPWR.t50 338.892
R2467 VPWR.n218 VPWR.n211 320.976
R2468 VPWR.n210 VPWR.n200 320.976
R2469 VPWR.n208 VPWR.n201 320.976
R2470 VPWR.n297 VPWR.n290 320.976
R2471 VPWR.n289 VPWR.n279 320.976
R2472 VPWR.n287 VPWR.n280 320.976
R2473 VPWR.n137 VPWR.n130 320.976
R2474 VPWR.n129 VPWR.n119 320.976
R2475 VPWR.n127 VPWR.n120 320.976
R2476 VPWR.n58 VPWR.n51 320.976
R2477 VPWR.n50 VPWR.n40 320.976
R2478 VPWR.n48 VPWR.n41 320.976
R2479 VPWR.n435 VPWR.n428 320.976
R2480 VPWR.n427 VPWR.n417 320.976
R2481 VPWR.n425 VPWR.n418 320.976
R2482 VPWR.n354 VPWR.n347 320.976
R2483 VPWR.n346 VPWR.n336 320.976
R2484 VPWR.n344 VPWR.n337 320.976
R2485 VPWR.n597 VPWR.n590 320.976
R2486 VPWR.n589 VPWR.n579 320.976
R2487 VPWR.n587 VPWR.n580 320.976
R2488 VPWR.n516 VPWR.n509 320.976
R2489 VPWR.n508 VPWR.n498 320.976
R2490 VPWR.n506 VPWR.n499 320.976
R2491 VPWR.n192 VPWR.t83 269.151
R2492 VPWR.n271 VPWR.t26 269.151
R2493 VPWR.n111 VPWR.t187 269.151
R2494 VPWR.n32 VPWR.t3 269.151
R2495 VPWR.n473 VPWR.t182 269.151
R2496 VPWR.n392 VPWR.t186 269.151
R2497 VPWR.n635 VPWR.t276 269.151
R2498 VPWR.n554 VPWR.t13 269.151
R2499 VPWR.n191 VPWR.t145 269.043
R2500 VPWR.n270 VPWR.t162 269.043
R2501 VPWR.n110 VPWR.t108 269.043
R2502 VPWR.n31 VPWR.t205 269.043
R2503 VPWR.n472 VPWR.t67 269.043
R2504 VPWR.n391 VPWR.t281 269.043
R2505 VPWR.n634 VPWR.t48 269.043
R2506 VPWR.n553 VPWR.t122 269.043
R2507 VPWR.n186 VPWR.t240 228.215
R2508 VPWR.n181 VPWR.t243 228.215
R2509 VPWR.n265 VPWR.t237 228.215
R2510 VPWR.n260 VPWR.t231 228.215
R2511 VPWR.n105 VPWR.t258 228.215
R2512 VPWR.n100 VPWR.t249 228.215
R2513 VPWR.n26 VPWR.t252 228.215
R2514 VPWR.n21 VPWR.t261 228.215
R2515 VPWR.n467 VPWR.t246 228.215
R2516 VPWR.n462 VPWR.t225 228.215
R2517 VPWR.n386 VPWR.t234 228.215
R2518 VPWR.n381 VPWR.t228 228.215
R2519 VPWR.n629 VPWR.t267 228.215
R2520 VPWR.n624 VPWR.t270 228.215
R2521 VPWR.n548 VPWR.t255 228.215
R2522 VPWR.n543 VPWR.t264 228.215
R2523 VPWR.t190 VPWR.n226 215.757
R2524 VPWR.n226 VPWR.t189 215.757
R2525 VPWR.t29 VPWR.n233 215.757
R2526 VPWR.n233 VPWR.t28 215.757
R2527 VPWR.t133 VPWR.n305 215.757
R2528 VPWR.n305 VPWR.t6 215.757
R2529 VPWR.t309 VPWR.n312 215.757
R2530 VPWR.n312 VPWR.t308 215.757
R2531 VPWR.t184 VPWR.n66 215.757
R2532 VPWR.n66 VPWR.t25 215.757
R2533 VPWR.t132 VPWR.n73 215.757
R2534 VPWR.n73 VPWR.t131 215.757
R2535 VPWR.t86 VPWR.n145 215.757
R2536 VPWR.n145 VPWR.t88 215.757
R2537 VPWR.t180 VPWR.n152 215.757
R2538 VPWR.n152 VPWR.t181 215.757
R2539 VPWR.t213 VPWR.n402 215.757
R2540 VPWR.n402 VPWR.t221 215.757
R2541 VPWR.t310 VPWR.n409 215.757
R2542 VPWR.n409 VPWR.t311 215.757
R2543 VPWR.t76 VPWR.n322 215.757
R2544 VPWR.n322 VPWR.t77 215.757
R2545 VPWR.t273 VPWR.n329 215.757
R2546 VPWR.n329 VPWR.t272 215.757
R2547 VPWR.t22 VPWR.n564 215.757
R2548 VPWR.n564 VPWR.t4 215.757
R2549 VPWR.t9 VPWR.n571 215.757
R2550 VPWR.n571 VPWR.t8 215.757
R2551 VPWR.t134 VPWR.n484 215.757
R2552 VPWR.n484 VPWR.t17 215.757
R2553 VPWR.t158 VPWR.n491 215.757
R2554 VPWR.n491 VPWR.t157 215.757
R2555 VPWR.n191 VPWR.t139 209.668
R2556 VPWR.n270 VPWR.t178 209.668
R2557 VPWR.n110 VPWR.t106 209.668
R2558 VPWR.n31 VPWR.t207 209.668
R2559 VPWR.n472 VPWR.t59 209.668
R2560 VPWR.n391 VPWR.t295 209.668
R2561 VPWR.n634 VPWR.t44 209.668
R2562 VPWR.n553 VPWR.t124 209.668
R2563 VPWR.n188 VPWR.n187 199.851
R2564 VPWR.n190 VPWR.n189 199.851
R2565 VPWR.n183 VPWR.n182 199.851
R2566 VPWR.n185 VPWR.n184 199.851
R2567 VPWR.n195 VPWR.n194 199.851
R2568 VPWR.n267 VPWR.n266 199.851
R2569 VPWR.n269 VPWR.n268 199.851
R2570 VPWR.n262 VPWR.n261 199.851
R2571 VPWR.n264 VPWR.n263 199.851
R2572 VPWR.n274 VPWR.n273 199.851
R2573 VPWR.n107 VPWR.n106 199.851
R2574 VPWR.n109 VPWR.n108 199.851
R2575 VPWR.n102 VPWR.n101 199.851
R2576 VPWR.n104 VPWR.n103 199.851
R2577 VPWR.n114 VPWR.n113 199.851
R2578 VPWR.n28 VPWR.n27 199.851
R2579 VPWR.n30 VPWR.n29 199.851
R2580 VPWR.n23 VPWR.n22 199.851
R2581 VPWR.n25 VPWR.n24 199.851
R2582 VPWR.n35 VPWR.n34 199.851
R2583 VPWR.n469 VPWR.n468 199.851
R2584 VPWR.n471 VPWR.n470 199.851
R2585 VPWR.n464 VPWR.n463 199.851
R2586 VPWR.n466 VPWR.n465 199.851
R2587 VPWR.n476 VPWR.n475 199.851
R2588 VPWR.n388 VPWR.n387 199.851
R2589 VPWR.n390 VPWR.n389 199.851
R2590 VPWR.n383 VPWR.n382 199.851
R2591 VPWR.n385 VPWR.n384 199.851
R2592 VPWR.n395 VPWR.n394 199.851
R2593 VPWR.n631 VPWR.n630 199.851
R2594 VPWR.n633 VPWR.n632 199.851
R2595 VPWR.n626 VPWR.n625 199.851
R2596 VPWR.n628 VPWR.n627 199.851
R2597 VPWR.n638 VPWR.n637 199.851
R2598 VPWR.n550 VPWR.n549 199.851
R2599 VPWR.n552 VPWR.n551 199.851
R2600 VPWR.n545 VPWR.n544 199.851
R2601 VPWR.n547 VPWR.n546 199.851
R2602 VPWR.n557 VPWR.n556 199.851
R2603 VPWR.n225 VPWR.n223 163.684
R2604 VPWR.n232 VPWR.n230 163.684
R2605 VPWR.n304 VPWR.n302 163.684
R2606 VPWR.n311 VPWR.n309 163.684
R2607 VPWR.n65 VPWR.n63 163.684
R2608 VPWR.n72 VPWR.n70 163.684
R2609 VPWR.n144 VPWR.n142 163.684
R2610 VPWR.n151 VPWR.n149 163.684
R2611 VPWR.n401 VPWR.n399 163.684
R2612 VPWR.n408 VPWR.n406 163.684
R2613 VPWR.n321 VPWR.n319 163.684
R2614 VPWR.n328 VPWR.n326 163.684
R2615 VPWR.n563 VPWR.n561 163.684
R2616 VPWR.n570 VPWR.n568 163.684
R2617 VPWR.n483 VPWR.n481 163.684
R2618 VPWR.n490 VPWR.n488 163.684
R2619 VPWR.n181 VPWR.t241 120.855
R2620 VPWR.n260 VPWR.t229 120.855
R2621 VPWR.n100 VPWR.t247 120.855
R2622 VPWR.n21 VPWR.t259 120.855
R2623 VPWR.n462 VPWR.t223 120.855
R2624 VPWR.n381 VPWR.t226 120.855
R2625 VPWR.n624 VPWR.t268 120.855
R2626 VPWR.n543 VPWR.t262 120.855
R2627 VPWR.n186 VPWR.t238 120.749
R2628 VPWR.n265 VPWR.t235 120.749
R2629 VPWR.n105 VPWR.t256 120.749
R2630 VPWR.n26 VPWR.t250 120.749
R2631 VPWR.n467 VPWR.t244 120.749
R2632 VPWR.n386 VPWR.t232 120.749
R2633 VPWR.n629 VPWR.t265 120.749
R2634 VPWR.n548 VPWR.t253 120.749
R2635 VPWR.n228 VPWR.n223 113.915
R2636 VPWR.n235 VPWR.n230 113.915
R2637 VPWR.n307 VPWR.n302 113.915
R2638 VPWR.n314 VPWR.n309 113.915
R2639 VPWR.n68 VPWR.n63 113.915
R2640 VPWR.n75 VPWR.n70 113.915
R2641 VPWR.n147 VPWR.n142 113.915
R2642 VPWR.n154 VPWR.n149 113.915
R2643 VPWR.n404 VPWR.n399 113.915
R2644 VPWR.n411 VPWR.n406 113.915
R2645 VPWR.n324 VPWR.n319 113.915
R2646 VPWR.n331 VPWR.n326 113.915
R2647 VPWR.n566 VPWR.n561 113.915
R2648 VPWR.n573 VPWR.n568 113.915
R2649 VPWR.n486 VPWR.n481 113.915
R2650 VPWR.n493 VPWR.n488 113.915
R2651 VPWR.n228 VPWR.n227 47.0382
R2652 VPWR.n235 VPWR.n234 47.0382
R2653 VPWR.n307 VPWR.n306 47.0382
R2654 VPWR.n314 VPWR.n313 47.0382
R2655 VPWR.n68 VPWR.n67 47.0382
R2656 VPWR.n75 VPWR.n74 47.0382
R2657 VPWR.n147 VPWR.n146 47.0382
R2658 VPWR.n154 VPWR.n153 47.0382
R2659 VPWR.n404 VPWR.n403 47.0382
R2660 VPWR.n411 VPWR.n410 47.0382
R2661 VPWR.n324 VPWR.n323 47.0382
R2662 VPWR.n331 VPWR.n330 47.0382
R2663 VPWR.n566 VPWR.n565 47.0382
R2664 VPWR.n573 VPWR.n572 47.0382
R2665 VPWR.n486 VPWR.n485 47.0382
R2666 VPWR.n493 VPWR.n492 47.0382
R2667 VPWR.n192 VPWR.n191 38.8096
R2668 VPWR.n271 VPWR.n270 38.8096
R2669 VPWR.n111 VPWR.n110 38.8096
R2670 VPWR.n32 VPWR.n31 38.8096
R2671 VPWR.n473 VPWR.n472 38.8096
R2672 VPWR.n392 VPWR.n391 38.8096
R2673 VPWR.n635 VPWR.n634 38.8096
R2674 VPWR.n554 VPWR.n553 38.8096
R2675 VPWR.n203 VPWR 35.5709
R2676 VPWR.n282 VPWR 35.5709
R2677 VPWR.n122 VPWR 35.5709
R2678 VPWR.n43 VPWR 35.5709
R2679 VPWR.n420 VPWR 35.5709
R2680 VPWR.n339 VPWR 35.5709
R2681 VPWR.n582 VPWR 35.5709
R2682 VPWR.n501 VPWR 35.5709
R2683 VPWR.n207 VPWR.n202 34.6358
R2684 VPWR.n220 VPWR.n219 34.6358
R2685 VPWR.n217 VPWR.n212 34.6358
R2686 VPWR.n286 VPWR.n281 34.6358
R2687 VPWR.n299 VPWR.n298 34.6358
R2688 VPWR.n296 VPWR.n291 34.6358
R2689 VPWR.n126 VPWR.n121 34.6358
R2690 VPWR.n139 VPWR.n138 34.6358
R2691 VPWR.n136 VPWR.n131 34.6358
R2692 VPWR.n47 VPWR.n42 34.6358
R2693 VPWR.n60 VPWR.n59 34.6358
R2694 VPWR.n57 VPWR.n52 34.6358
R2695 VPWR.n424 VPWR.n419 34.6358
R2696 VPWR.n437 VPWR.n436 34.6358
R2697 VPWR.n434 VPWR.n429 34.6358
R2698 VPWR.n343 VPWR.n338 34.6358
R2699 VPWR.n356 VPWR.n355 34.6358
R2700 VPWR.n353 VPWR.n348 34.6358
R2701 VPWR.n586 VPWR.n581 34.6358
R2702 VPWR.n599 VPWR.n598 34.6358
R2703 VPWR.n596 VPWR.n591 34.6358
R2704 VPWR.n505 VPWR.n500 34.6358
R2705 VPWR.n518 VPWR.n517 34.6358
R2706 VPWR.n515 VPWR.n510 34.6358
R2707 VPWR.n210 VPWR.n209 32.0005
R2708 VPWR.n289 VPWR.n288 32.0005
R2709 VPWR.n129 VPWR.n128 32.0005
R2710 VPWR.n50 VPWR.n49 32.0005
R2711 VPWR.n427 VPWR.n426 32.0005
R2712 VPWR.n346 VPWR.n345 32.0005
R2713 VPWR.n589 VPWR.n588 32.0005
R2714 VPWR.n508 VPWR.n507 32.0005
R2715 VPWR.n209 VPWR.n208 31.2476
R2716 VPWR.n288 VPWR.n287 31.2476
R2717 VPWR.n128 VPWR.n127 31.2476
R2718 VPWR.n49 VPWR.n48 31.2476
R2719 VPWR.n426 VPWR.n425 31.2476
R2720 VPWR.n345 VPWR.n344 31.2476
R2721 VPWR.n588 VPWR.n587 31.2476
R2722 VPWR.n507 VPWR.n506 31.2476
R2723 VPWR.n187 VPWR.t138 28.5655
R2724 VPWR.n187 VPWR.t156 28.5655
R2725 VPWR.n189 VPWR.t148 28.5655
R2726 VPWR.n189 VPWR.t152 28.5655
R2727 VPWR.n182 VPWR.t144 28.5655
R2728 VPWR.n182 VPWR.t150 28.5655
R2729 VPWR.n184 VPWR.t154 28.5655
R2730 VPWR.n184 VPWR.t142 28.5655
R2731 VPWR.n194 VPWR.t140 28.5655
R2732 VPWR.n194 VPWR.t146 28.5655
R2733 VPWR.n266 VPWR.t171 28.5655
R2734 VPWR.n266 VPWR.t177 28.5655
R2735 VPWR.n268 VPWR.t167 28.5655
R2736 VPWR.n268 VPWR.t173 28.5655
R2737 VPWR.n261 VPWR.t165 28.5655
R2738 VPWR.n261 VPWR.t169 28.5655
R2739 VPWR.n263 VPWR.t175 28.5655
R2740 VPWR.n263 VPWR.t161 28.5655
R2741 VPWR.n273 VPWR.t179 28.5655
R2742 VPWR.n273 VPWR.t163 28.5655
R2743 VPWR.n106 VPWR.t97 28.5655
R2744 VPWR.n106 VPWR.t105 28.5655
R2745 VPWR.n108 VPWR.t91 28.5655
R2746 VPWR.n108 VPWR.t99 28.5655
R2747 VPWR.n101 VPWR.t93 28.5655
R2748 VPWR.n101 VPWR.t95 28.5655
R2749 VPWR.n103 VPWR.t103 28.5655
R2750 VPWR.n103 VPWR.t101 28.5655
R2751 VPWR.n113 VPWR.t107 28.5655
R2752 VPWR.n113 VPWR.t109 28.5655
R2753 VPWR.n27 VPWR.t200 28.5655
R2754 VPWR.n27 VPWR.t204 28.5655
R2755 VPWR.n29 VPWR.t212 28.5655
R2756 VPWR.n29 VPWR.t196 28.5655
R2757 VPWR.n22 VPWR.t210 28.5655
R2758 VPWR.n22 VPWR.t194 28.5655
R2759 VPWR.n24 VPWR.t198 28.5655
R2760 VPWR.n24 VPWR.t202 28.5655
R2761 VPWR.n34 VPWR.t208 28.5655
R2762 VPWR.n34 VPWR.t206 28.5655
R2763 VPWR.n468 VPWR.t58 28.5655
R2764 VPWR.n468 VPWR.t56 28.5655
R2765 VPWR.n470 VPWR.t64 28.5655
R2766 VPWR.n470 VPWR.t72 28.5655
R2767 VPWR.n463 VPWR.t66 28.5655
R2768 VPWR.n463 VPWR.t70 28.5655
R2769 VPWR.n465 VPWR.t74 28.5655
R2770 VPWR.n465 VPWR.t62 28.5655
R2771 VPWR.n475 VPWR.t60 28.5655
R2772 VPWR.n475 VPWR.t68 28.5655
R2773 VPWR.n387 VPWR.t292 28.5655
R2774 VPWR.n387 VPWR.t294 28.5655
R2775 VPWR.n389 VPWR.t280 28.5655
R2776 VPWR.n389 VPWR.t288 28.5655
R2777 VPWR.n382 VPWR.t286 28.5655
R2778 VPWR.n382 VPWR.t284 28.5655
R2779 VPWR.n384 VPWR.t290 28.5655
R2780 VPWR.n384 VPWR.t278 28.5655
R2781 VPWR.n394 VPWR.t296 28.5655
R2782 VPWR.n394 VPWR.t282 28.5655
R2783 VPWR.n630 VPWR.t39 28.5655
R2784 VPWR.n630 VPWR.t43 28.5655
R2785 VPWR.n632 VPWR.t33 28.5655
R2786 VPWR.n632 VPWR.t31 28.5655
R2787 VPWR.n625 VPWR.t47 28.5655
R2788 VPWR.n625 VPWR.t37 28.5655
R2789 VPWR.n627 VPWR.t35 28.5655
R2790 VPWR.n627 VPWR.t41 28.5655
R2791 VPWR.n637 VPWR.t45 28.5655
R2792 VPWR.n637 VPWR.t49 28.5655
R2793 VPWR.n549 VPWR.t117 28.5655
R2794 VPWR.n549 VPWR.t121 28.5655
R2795 VPWR.n551 VPWR.t111 28.5655
R2796 VPWR.n551 VPWR.t129 28.5655
R2797 VPWR.n544 VPWR.t127 28.5655
R2798 VPWR.n544 VPWR.t113 28.5655
R2799 VPWR.n546 VPWR.t115 28.5655
R2800 VPWR.n546 VPWR.t119 28.5655
R2801 VPWR.n556 VPWR.t125 28.5655
R2802 VPWR.n556 VPWR.t123 28.5655
R2803 VPWR.n211 VPWR.t53 26.5955
R2804 VPWR.n211 VPWR.t89 26.5955
R2805 VPWR.n200 VPWR.t303 26.5955
R2806 VPWR.n200 VPWR.t0 26.5955
R2807 VPWR.n201 VPWR.t12 26.5955
R2808 VPWR.n201 VPWR.t85 26.5955
R2809 VPWR.n290 VPWR.t275 26.5955
R2810 VPWR.n290 VPWR.t81 26.5955
R2811 VPWR.n279 VPWR.t188 26.5955
R2812 VPWR.n279 VPWR.t14 26.5955
R2813 VPWR.n280 VPWR.t274 26.5955
R2814 VPWR.n280 VPWR.t298 26.5955
R2815 VPWR.n130 VPWR.t21 26.5955
R2816 VPWR.n130 VPWR.t5 26.5955
R2817 VPWR.n119 VPWR.t159 26.5955
R2818 VPWR.n119 VPWR.t80 26.5955
R2819 VPWR.n120 VPWR.t52 26.5955
R2820 VPWR.n120 VPWR.t54 26.5955
R2821 VPWR.n51 VPWR.t136 26.5955
R2822 VPWR.n51 VPWR.t20 26.5955
R2823 VPWR.n40 VPWR.t84 26.5955
R2824 VPWR.n40 VPWR.t79 26.5955
R2825 VPWR.n41 VPWR.t305 26.5955
R2826 VPWR.n41 VPWR.t87 26.5955
R2827 VPWR.n428 VPWR.t220 26.5955
R2828 VPWR.n428 VPWR.t222 26.5955
R2829 VPWR.n417 VPWR.t219 26.5955
R2830 VPWR.n417 VPWR.t217 26.5955
R2831 VPWR.n418 VPWR.t216 26.5955
R2832 VPWR.n418 VPWR.t214 26.5955
R2833 VPWR.n347 VPWR.t75 26.5955
R2834 VPWR.n347 VPWR.t19 26.5955
R2835 VPWR.n336 VPWR.t135 26.5955
R2836 VPWR.n336 VPWR.t18 26.5955
R2837 VPWR.n337 VPWR.t78 26.5955
R2838 VPWR.n337 VPWR.t304 26.5955
R2839 VPWR.n590 VPWR.t271 26.5955
R2840 VPWR.n590 VPWR.t2 26.5955
R2841 VPWR.n579 VPWR.t23 26.5955
R2842 VPWR.n579 VPWR.t297 26.5955
R2843 VPWR.n580 VPWR.t10 26.5955
R2844 VPWR.n580 VPWR.t11 26.5955
R2845 VPWR.n509 VPWR.t300 26.5955
R2846 VPWR.n509 VPWR.t7 26.5955
R2847 VPWR.n498 VPWR.t16 26.5955
R2848 VPWR.n498 VPWR.t302 26.5955
R2849 VPWR.n499 VPWR.t299 26.5955
R2850 VPWR.n499 VPWR.t191 26.5955
R2851 VPWR.n219 VPWR.n218 25.977
R2852 VPWR.n298 VPWR.n297 25.977
R2853 VPWR.n138 VPWR.n137 25.977
R2854 VPWR.n59 VPWR.n58 25.977
R2855 VPWR.n436 VPWR.n435 25.977
R2856 VPWR.n355 VPWR.n354 25.977
R2857 VPWR.n598 VPWR.n597 25.977
R2858 VPWR.n517 VPWR.n516 25.977
R2859 VPWR.n226 VPWR.n224 20.5561
R2860 VPWR.n233 VPWR.n231 20.5561
R2861 VPWR.n305 VPWR.n303 20.5561
R2862 VPWR.n312 VPWR.n310 20.5561
R2863 VPWR.n66 VPWR.n64 20.5561
R2864 VPWR.n73 VPWR.n71 20.5561
R2865 VPWR.n145 VPWR.n143 20.5561
R2866 VPWR.n152 VPWR.n150 20.5561
R2867 VPWR.n402 VPWR.n400 20.5561
R2868 VPWR.n409 VPWR.n407 20.5561
R2869 VPWR.n322 VPWR.n320 20.5561
R2870 VPWR.n329 VPWR.n327 20.5561
R2871 VPWR.n564 VPWR.n562 20.5561
R2872 VPWR.n571 VPWR.n569 20.5561
R2873 VPWR.n484 VPWR.n482 20.5561
R2874 VPWR.n491 VPWR.n489 20.5561
R2875 VPWR.n203 VPWR.n202 18.824
R2876 VPWR.n282 VPWR.n281 18.824
R2877 VPWR.n122 VPWR.n121 18.824
R2878 VPWR.n43 VPWR.n42 18.824
R2879 VPWR.n420 VPWR.n419 18.824
R2880 VPWR.n339 VPWR.n338 18.824
R2881 VPWR.n582 VPWR.n581 18.824
R2882 VPWR.n501 VPWR.n500 18.824
R2883 VPWR.n224 VPWR.n223 18.7435
R2884 VPWR.n231 VPWR.n230 18.7435
R2885 VPWR.n303 VPWR.n302 18.7435
R2886 VPWR.n310 VPWR.n309 18.7435
R2887 VPWR.n64 VPWR.n63 18.7435
R2888 VPWR.n71 VPWR.n70 18.7435
R2889 VPWR.n143 VPWR.n142 18.7435
R2890 VPWR.n150 VPWR.n149 18.7435
R2891 VPWR.n400 VPWR.n399 18.7435
R2892 VPWR.n407 VPWR.n406 18.7435
R2893 VPWR.n320 VPWR.n319 18.7435
R2894 VPWR.n327 VPWR.n326 18.7435
R2895 VPWR.n562 VPWR.n561 18.7435
R2896 VPWR.n569 VPWR.n568 18.7435
R2897 VPWR.n482 VPWR.n481 18.7435
R2898 VPWR.n489 VPWR.n488 18.7435
R2899 VPWR.n213 VPWR.n212 13.5534
R2900 VPWR.n292 VPWR.n291 13.5534
R2901 VPWR.n132 VPWR.n131 13.5534
R2902 VPWR.n53 VPWR.n52 13.5534
R2903 VPWR.n430 VPWR.n429 13.5534
R2904 VPWR.n349 VPWR.n348 13.5534
R2905 VPWR.n592 VPWR.n591 13.5534
R2906 VPWR.n511 VPWR.n510 13.5534
R2907 VPWR VPWR.n228 11.4981
R2908 VPWR VPWR.n235 11.4981
R2909 VPWR VPWR.n307 11.4981
R2910 VPWR VPWR.n314 11.4981
R2911 VPWR VPWR.n68 11.4981
R2912 VPWR VPWR.n75 11.4981
R2913 VPWR VPWR.n147 11.4981
R2914 VPWR VPWR.n154 11.4981
R2915 VPWR VPWR.n404 11.4981
R2916 VPWR VPWR.n411 11.4981
R2917 VPWR VPWR.n324 11.4981
R2918 VPWR VPWR.n331 11.4981
R2919 VPWR VPWR.n566 11.4981
R2920 VPWR VPWR.n573 11.4981
R2921 VPWR VPWR.n486 11.4981
R2922 VPWR VPWR.n493 11.4981
R2923 VPWR.n214 VPWR.n213 11.1829
R2924 VPWR.n293 VPWR.n292 11.1829
R2925 VPWR.n133 VPWR.n132 11.1829
R2926 VPWR.n54 VPWR.n53 11.1829
R2927 VPWR.n431 VPWR.n430 11.1829
R2928 VPWR.n350 VPWR.n349 11.1829
R2929 VPWR.n593 VPWR.n592 11.1829
R2930 VPWR.n512 VPWR.n511 11.1829
R2931 VPWR.n204 VPWR.n203 9.3005
R2932 VPWR.n205 VPWR.n202 9.3005
R2933 VPWR.n207 VPWR.n206 9.3005
R2934 VPWR.n209 VPWR.n198 9.3005
R2935 VPWR.n221 VPWR.n220 9.3005
R2936 VPWR.n219 VPWR.n199 9.3005
R2937 VPWR.n217 VPWR.n216 9.3005
R2938 VPWR.n215 VPWR.n212 9.3005
R2939 VPWR.n283 VPWR.n282 9.3005
R2940 VPWR.n284 VPWR.n281 9.3005
R2941 VPWR.n286 VPWR.n285 9.3005
R2942 VPWR.n288 VPWR.n277 9.3005
R2943 VPWR.n300 VPWR.n299 9.3005
R2944 VPWR.n298 VPWR.n278 9.3005
R2945 VPWR.n296 VPWR.n295 9.3005
R2946 VPWR.n294 VPWR.n291 9.3005
R2947 VPWR.n123 VPWR.n122 9.3005
R2948 VPWR.n124 VPWR.n121 9.3005
R2949 VPWR.n126 VPWR.n125 9.3005
R2950 VPWR.n128 VPWR.n117 9.3005
R2951 VPWR.n140 VPWR.n139 9.3005
R2952 VPWR.n138 VPWR.n118 9.3005
R2953 VPWR.n136 VPWR.n135 9.3005
R2954 VPWR.n134 VPWR.n131 9.3005
R2955 VPWR.n44 VPWR.n43 9.3005
R2956 VPWR.n45 VPWR.n42 9.3005
R2957 VPWR.n47 VPWR.n46 9.3005
R2958 VPWR.n49 VPWR.n38 9.3005
R2959 VPWR.n61 VPWR.n60 9.3005
R2960 VPWR.n59 VPWR.n39 9.3005
R2961 VPWR.n57 VPWR.n56 9.3005
R2962 VPWR.n55 VPWR.n52 9.3005
R2963 VPWR.n421 VPWR.n420 9.3005
R2964 VPWR.n422 VPWR.n419 9.3005
R2965 VPWR.n424 VPWR.n423 9.3005
R2966 VPWR.n426 VPWR.n415 9.3005
R2967 VPWR.n438 VPWR.n437 9.3005
R2968 VPWR.n436 VPWR.n416 9.3005
R2969 VPWR.n434 VPWR.n433 9.3005
R2970 VPWR.n432 VPWR.n429 9.3005
R2971 VPWR.n340 VPWR.n339 9.3005
R2972 VPWR.n341 VPWR.n338 9.3005
R2973 VPWR.n343 VPWR.n342 9.3005
R2974 VPWR.n345 VPWR.n334 9.3005
R2975 VPWR.n357 VPWR.n356 9.3005
R2976 VPWR.n355 VPWR.n335 9.3005
R2977 VPWR.n353 VPWR.n352 9.3005
R2978 VPWR.n351 VPWR.n348 9.3005
R2979 VPWR.n583 VPWR.n582 9.3005
R2980 VPWR.n584 VPWR.n581 9.3005
R2981 VPWR.n586 VPWR.n585 9.3005
R2982 VPWR.n588 VPWR.n577 9.3005
R2983 VPWR.n600 VPWR.n599 9.3005
R2984 VPWR.n598 VPWR.n578 9.3005
R2985 VPWR.n596 VPWR.n595 9.3005
R2986 VPWR.n594 VPWR.n591 9.3005
R2987 VPWR.n502 VPWR.n501 9.3005
R2988 VPWR.n503 VPWR.n500 9.3005
R2989 VPWR.n505 VPWR.n504 9.3005
R2990 VPWR.n507 VPWR.n496 9.3005
R2991 VPWR.n519 VPWR.n518 9.3005
R2992 VPWR.n517 VPWR.n497 9.3005
R2993 VPWR.n515 VPWR.n514 9.3005
R2994 VPWR.n513 VPWR.n510 9.3005
R2995 VPWR.n218 VPWR.n217 8.65932
R2996 VPWR.n297 VPWR.n296 8.65932
R2997 VPWR.n137 VPWR.n136 8.65932
R2998 VPWR.n58 VPWR.n57 8.65932
R2999 VPWR.n435 VPWR.n434 8.65932
R3000 VPWR.n354 VPWR.n353 8.65932
R3001 VPWR.n597 VPWR.n596 8.65932
R3002 VPWR.n516 VPWR.n515 8.65932
R3003 VPWR.n78 VPWR 5.89271
R3004 VPWR.n168 VPWR.n165 5.0005
R3005 VPWR.n174 VPWR.n165 5.0005
R3006 VPWR.n247 VPWR.n244 5.0005
R3007 VPWR.n253 VPWR.n244 5.0005
R3008 VPWR.n87 VPWR.n84 5.0005
R3009 VPWR.n93 VPWR.n84 5.0005
R3010 VPWR.n8 VPWR.n5 5.0005
R3011 VPWR.n14 VPWR.n5 5.0005
R3012 VPWR.n449 VPWR.n446 5.0005
R3013 VPWR.n455 VPWR.n446 5.0005
R3014 VPWR.n368 VPWR.n365 5.0005
R3015 VPWR.n374 VPWR.n365 5.0005
R3016 VPWR.n611 VPWR.n608 5.0005
R3017 VPWR.n617 VPWR.n608 5.0005
R3018 VPWR.n530 VPWR.n527 5.0005
R3019 VPWR.n536 VPWR.n527 5.0005
R3020 VPWR.n159 VPWR 4.95117
R3021 VPWR.n167 VPWR.n164 4.86892
R3022 VPWR.n166 VPWR.n164 4.86892
R3023 VPWR.n246 VPWR.n243 4.86892
R3024 VPWR.n245 VPWR.n243 4.86892
R3025 VPWR.n86 VPWR.n83 4.86892
R3026 VPWR.n85 VPWR.n83 4.86892
R3027 VPWR.n7 VPWR.n4 4.86892
R3028 VPWR.n6 VPWR.n4 4.86892
R3029 VPWR.n448 VPWR.n445 4.86892
R3030 VPWR.n447 VPWR.n445 4.86892
R3031 VPWR.n367 VPWR.n364 4.86892
R3032 VPWR.n366 VPWR.n364 4.86892
R3033 VPWR.n610 VPWR.n607 4.86892
R3034 VPWR.n609 VPWR.n607 4.86892
R3035 VPWR.n529 VPWR.n526 4.86892
R3036 VPWR.n528 VPWR.n526 4.86892
R3037 VPWR.n480 VPWR 3.8545
R3038 VPWR.n208 VPWR.n207 3.38874
R3039 VPWR.n287 VPWR.n286 3.38874
R3040 VPWR.n127 VPWR.n126 3.38874
R3041 VPWR.n48 VPWR.n47 3.38874
R3042 VPWR.n425 VPWR.n424 3.38874
R3043 VPWR.n344 VPWR.n343 3.38874
R3044 VPWR.n587 VPWR.n586 3.38874
R3045 VPWR.n506 VPWR.n505 3.38874
R3046 VPWR.n237 VPWR.n236 3.28283
R3047 VPWR.n316 VPWR.n315 3.28283
R3048 VPWR.n77 VPWR.n76 3.28283
R3049 VPWR.n156 VPWR.n155 3.28283
R3050 VPWR.n413 VPWR.n412 3.28283
R3051 VPWR.n333 VPWR.n332 3.28283
R3052 VPWR.n575 VPWR.n574 3.28283
R3053 VPWR.n495 VPWR.n494 3.28283
R3054 VPWR.n237 VPWR.n229 3.19667
R3055 VPWR.n316 VPWR.n308 3.19667
R3056 VPWR.n77 VPWR.n69 3.19667
R3057 VPWR.n156 VPWR.n148 3.19667
R3058 VPWR.n413 VPWR.n405 3.19667
R3059 VPWR.n333 VPWR.n325 3.19667
R3060 VPWR.n575 VPWR.n567 3.19667
R3061 VPWR.n495 VPWR.n487 3.19667
R3062 VPWR.n642 VPWR 2.7265
R3063 VPWR.n220 VPWR.n210 2.63579
R3064 VPWR.n299 VPWR.n289 2.63579
R3065 VPWR.n139 VPWR.n129 2.63579
R3066 VPWR.n60 VPWR.n50 2.63579
R3067 VPWR.n437 VPWR.n427 2.63579
R3068 VPWR.n356 VPWR.n346 2.63579
R3069 VPWR.n599 VPWR.n589 2.63579
R3070 VPWR.n518 VPWR.n508 2.63579
R3071 VPWR.n642 VPWR 2.5385
R3072 VPWR.n179 VPWR.n161 2.4755
R3073 VPWR.n169 VPWR.n161 2.4755
R3074 VPWR.n258 VPWR.n240 2.4755
R3075 VPWR.n248 VPWR.n240 2.4755
R3076 VPWR.n98 VPWR.n80 2.4755
R3077 VPWR.n88 VPWR.n80 2.4755
R3078 VPWR.n19 VPWR.n1 2.4755
R3079 VPWR.n9 VPWR.n1 2.4755
R3080 VPWR.n460 VPWR.n442 2.4755
R3081 VPWR.n450 VPWR.n442 2.4755
R3082 VPWR.n379 VPWR.n361 2.4755
R3083 VPWR.n369 VPWR.n361 2.4755
R3084 VPWR.n622 VPWR.n604 2.4755
R3085 VPWR.n612 VPWR.n604 2.4755
R3086 VPWR.n541 VPWR.n523 2.4755
R3087 VPWR.n531 VPWR.n523 2.4755
R3088 VPWR.n169 VPWR.n160 2.463
R3089 VPWR.n248 VPWR.n239 2.463
R3090 VPWR.n88 VPWR.n79 2.463
R3091 VPWR.n9 VPWR.n0 2.463
R3092 VPWR.n450 VPWR.n441 2.463
R3093 VPWR.n369 VPWR.n360 2.463
R3094 VPWR.n612 VPWR.n603 2.463
R3095 VPWR.n531 VPWR.n522 2.463
R3096 VPWR.n177 VPWR.n176 2.34227
R3097 VPWR.n176 VPWR.n175 2.34227
R3098 VPWR.n172 VPWR.n171 2.34227
R3099 VPWR.n173 VPWR.n172 2.34227
R3100 VPWR.n256 VPWR.n255 2.34227
R3101 VPWR.n255 VPWR.n254 2.34227
R3102 VPWR.n251 VPWR.n250 2.34227
R3103 VPWR.n252 VPWR.n251 2.34227
R3104 VPWR.n96 VPWR.n95 2.34227
R3105 VPWR.n95 VPWR.n94 2.34227
R3106 VPWR.n91 VPWR.n90 2.34227
R3107 VPWR.n92 VPWR.n91 2.34227
R3108 VPWR.n17 VPWR.n16 2.34227
R3109 VPWR.n16 VPWR.n15 2.34227
R3110 VPWR.n12 VPWR.n11 2.34227
R3111 VPWR.n13 VPWR.n12 2.34227
R3112 VPWR.n458 VPWR.n457 2.34227
R3113 VPWR.n457 VPWR.n456 2.34227
R3114 VPWR.n453 VPWR.n452 2.34227
R3115 VPWR.n454 VPWR.n453 2.34227
R3116 VPWR.n377 VPWR.n376 2.34227
R3117 VPWR.n376 VPWR.n375 2.34227
R3118 VPWR.n372 VPWR.n371 2.34227
R3119 VPWR.n373 VPWR.n372 2.34227
R3120 VPWR.n620 VPWR.n619 2.34227
R3121 VPWR.n619 VPWR.n618 2.34227
R3122 VPWR.n615 VPWR.n614 2.34227
R3123 VPWR.n616 VPWR.n615 2.34227
R3124 VPWR.n539 VPWR.n538 2.34227
R3125 VPWR.n538 VPWR.n537 2.34227
R3126 VPWR.n534 VPWR.n533 2.34227
R3127 VPWR.n535 VPWR.n534 2.34227
R3128 VPWR.n180 VPWR.n160 2.10363
R3129 VPWR.n259 VPWR.n239 2.10363
R3130 VPWR.n99 VPWR.n79 2.10363
R3131 VPWR.n20 VPWR.n0 2.10363
R3132 VPWR.n461 VPWR.n441 2.10363
R3133 VPWR.n380 VPWR.n360 2.10363
R3134 VPWR.n623 VPWR.n603 2.10363
R3135 VPWR.n542 VPWR.n522 2.10363
R3136 VPWR.n178 VPWR.n177 1.93989
R3137 VPWR.n257 VPWR.n256 1.93989
R3138 VPWR.n97 VPWR.n96 1.93989
R3139 VPWR.n18 VPWR.n17 1.93989
R3140 VPWR.n459 VPWR.n458 1.93989
R3141 VPWR.n378 VPWR.n377 1.93989
R3142 VPWR.n621 VPWR.n620 1.93989
R3143 VPWR.n540 VPWR.n539 1.93989
R3144 VPWR.n238 VPWR.n222 1.02714
R3145 VPWR.n317 VPWR.n301 1.02714
R3146 VPWR.n157 VPWR.n141 1.02714
R3147 VPWR.n78 VPWR.n62 1.02714
R3148 VPWR.n440 VPWR.n439 1.02714
R3149 VPWR.n359 VPWR.n358 1.02714
R3150 VPWR.n602 VPWR.n601 1.02714
R3151 VPWR.n521 VPWR.n520 1.02714
R3152 VPWR.n167 VPWR.n162 0.970197
R3153 VPWR.n171 VPWR.n170 0.970197
R3154 VPWR.n168 VPWR.n163 0.970197
R3155 VPWR.n246 VPWR.n241 0.970197
R3156 VPWR.n250 VPWR.n249 0.970197
R3157 VPWR.n247 VPWR.n242 0.970197
R3158 VPWR.n86 VPWR.n81 0.970197
R3159 VPWR.n90 VPWR.n89 0.970197
R3160 VPWR.n87 VPWR.n82 0.970197
R3161 VPWR.n7 VPWR.n2 0.970197
R3162 VPWR.n11 VPWR.n10 0.970197
R3163 VPWR.n8 VPWR.n3 0.970197
R3164 VPWR.n448 VPWR.n443 0.970197
R3165 VPWR.n452 VPWR.n451 0.970197
R3166 VPWR.n449 VPWR.n444 0.970197
R3167 VPWR.n367 VPWR.n362 0.970197
R3168 VPWR.n371 VPWR.n370 0.970197
R3169 VPWR.n368 VPWR.n363 0.970197
R3170 VPWR.n610 VPWR.n605 0.970197
R3171 VPWR.n614 VPWR.n613 0.970197
R3172 VPWR.n611 VPWR.n606 0.970197
R3173 VPWR.n529 VPWR.n524 0.970197
R3174 VPWR.n533 VPWR.n532 0.970197
R3175 VPWR.n530 VPWR.n525 0.970197
R3176 VPWR.n183 VPWR.n181 0.890989
R3177 VPWR.n262 VPWR.n260 0.890989
R3178 VPWR.n102 VPWR.n100 0.890989
R3179 VPWR.n23 VPWR.n21 0.890989
R3180 VPWR.n464 VPWR.n462 0.890989
R3181 VPWR.n383 VPWR.n381 0.890989
R3182 VPWR.n626 VPWR.n624 0.890989
R3183 VPWR.n545 VPWR.n543 0.890989
R3184 VPWR.n642 VPWR.n480 0.877833
R3185 VPWR.n480 VPWR.n318 0.8465
R3186 VPWR.n188 VPWR.n186 0.760446
R3187 VPWR.n267 VPWR.n265 0.760446
R3188 VPWR.n107 VPWR.n105 0.760446
R3189 VPWR.n28 VPWR.n26 0.760446
R3190 VPWR.n469 VPWR.n467 0.760446
R3191 VPWR.n388 VPWR.n386 0.760446
R3192 VPWR.n631 VPWR.n629 0.760446
R3193 VPWR.n550 VPWR.n548 0.760446
R3194 VPWR.n159 VPWR.n158 0.689833
R3195 VPWR.n190 VPWR.n188 0.40675
R3196 VPWR.n185 VPWR.n183 0.40675
R3197 VPWR.n195 VPWR.n185 0.40675
R3198 VPWR.n269 VPWR.n267 0.40675
R3199 VPWR.n264 VPWR.n262 0.40675
R3200 VPWR.n274 VPWR.n264 0.40675
R3201 VPWR.n109 VPWR.n107 0.40675
R3202 VPWR.n104 VPWR.n102 0.40675
R3203 VPWR.n114 VPWR.n104 0.40675
R3204 VPWR.n30 VPWR.n28 0.40675
R3205 VPWR.n25 VPWR.n23 0.40675
R3206 VPWR.n35 VPWR.n25 0.40675
R3207 VPWR.n471 VPWR.n469 0.40675
R3208 VPWR.n466 VPWR.n464 0.40675
R3209 VPWR.n476 VPWR.n466 0.40675
R3210 VPWR.n390 VPWR.n388 0.40675
R3211 VPWR.n385 VPWR.n383 0.40675
R3212 VPWR.n395 VPWR.n385 0.40675
R3213 VPWR.n633 VPWR.n631 0.40675
R3214 VPWR.n628 VPWR.n626 0.40675
R3215 VPWR.n638 VPWR.n628 0.40675
R3216 VPWR.n552 VPWR.n550 0.40675
R3217 VPWR.n547 VPWR.n545 0.40675
R3218 VPWR.n557 VPWR.n547 0.40675
R3219 VPWR.n521 VPWR.n495 0.397508
R3220 VPWR.n359 VPWR.n333 0.383506
R3221 VPWR.n180 VPWR.n179 0.359875
R3222 VPWR.n259 VPWR.n258 0.359875
R3223 VPWR.n99 VPWR.n98 0.359875
R3224 VPWR.n20 VPWR.n19 0.359875
R3225 VPWR.n461 VPWR.n460 0.359875
R3226 VPWR.n380 VPWR.n379 0.359875
R3227 VPWR.n623 VPWR.n622 0.359875
R3228 VPWR.n542 VPWR.n541 0.359875
R3229 VPWR.n157 VPWR.n156 0.3415
R3230 VPWR.n78 VPWR.n77 0.3415
R3231 VPWR.n317 VPWR.n316 0.3415
R3232 VPWR.n238 VPWR.n237 0.3415
R3233 VPWR.n414 VPWR.n413 0.3415
R3234 VPWR.n576 VPWR.n575 0.3415
R3235 VPWR.n163 VPWR.n161 0.258833
R3236 VPWR.n162 VPWR.n160 0.258833
R3237 VPWR.n242 VPWR.n240 0.258833
R3238 VPWR.n241 VPWR.n239 0.258833
R3239 VPWR.n82 VPWR.n80 0.258833
R3240 VPWR.n81 VPWR.n79 0.258833
R3241 VPWR.n3 VPWR.n1 0.258833
R3242 VPWR.n2 VPWR.n0 0.258833
R3243 VPWR.n444 VPWR.n442 0.258833
R3244 VPWR.n443 VPWR.n441 0.258833
R3245 VPWR.n363 VPWR.n361 0.258833
R3246 VPWR.n362 VPWR.n360 0.258833
R3247 VPWR.n606 VPWR.n604 0.258833
R3248 VPWR.n605 VPWR.n603 0.258833
R3249 VPWR.n525 VPWR.n523 0.258833
R3250 VPWR.n524 VPWR.n522 0.258833
R3251 VPWR.n195 VPWR.n193 0.208833
R3252 VPWR.n274 VPWR.n272 0.208833
R3253 VPWR.n114 VPWR.n112 0.208833
R3254 VPWR.n35 VPWR.n33 0.208833
R3255 VPWR.n476 VPWR.n474 0.208833
R3256 VPWR.n395 VPWR.n393 0.208833
R3257 VPWR.n638 VPWR.n636 0.208833
R3258 VPWR.n557 VPWR.n555 0.208833
R3259 VPWR.n193 VPWR.n190 0.188
R3260 VPWR.n272 VPWR.n269 0.188
R3261 VPWR.n112 VPWR.n109 0.188
R3262 VPWR.n33 VPWR.n30 0.188
R3263 VPWR.n474 VPWR.n471 0.188
R3264 VPWR.n393 VPWR.n390 0.188
R3265 VPWR.n636 VPWR.n633 0.188
R3266 VPWR.n555 VPWR.n552 0.188
R3267 VPWR.n193 VPWR.n192 0.1865
R3268 VPWR.n272 VPWR.n271 0.1865
R3269 VPWR.n112 VPWR.n111 0.1865
R3270 VPWR.n33 VPWR.n32 0.1865
R3271 VPWR.n474 VPWR.n473 0.1865
R3272 VPWR.n393 VPWR.n392 0.1865
R3273 VPWR.n636 VPWR.n635 0.1865
R3274 VPWR.n555 VPWR.n554 0.1865
R3275 VPWR.n560 VPWR.n521 0.184975
R3276 VPWR.n641 VPWR.n602 0.184975
R3277 VPWR.n642 VPWR 0.178395
R3278 VPWR.n576 VPWR 0.167428
R3279 VPWR.n398 VPWR.n359 0.138856
R3280 VPWR.n479 VPWR.n440 0.138856
R3281 VPWR.n480 VPWR 0.137564
R3282 VPWR.n170 VPWR.n169 0.121279
R3283 VPWR.n179 VPWR.n178 0.121279
R3284 VPWR.n249 VPWR.n248 0.121279
R3285 VPWR.n258 VPWR.n257 0.121279
R3286 VPWR.n89 VPWR.n88 0.121279
R3287 VPWR.n98 VPWR.n97 0.121279
R3288 VPWR.n10 VPWR.n9 0.121279
R3289 VPWR.n19 VPWR.n18 0.121279
R3290 VPWR.n451 VPWR.n450 0.121279
R3291 VPWR.n460 VPWR.n459 0.121279
R3292 VPWR.n370 VPWR.n369 0.121279
R3293 VPWR.n379 VPWR.n378 0.121279
R3294 VPWR.n613 VPWR.n612 0.121279
R3295 VPWR.n622 VPWR.n621 0.121279
R3296 VPWR.n532 VPWR.n531 0.121279
R3297 VPWR.n541 VPWR.n540 0.121279
R3298 VPWR.n205 VPWR.n204 0.120292
R3299 VPWR.n206 VPWR.n205 0.120292
R3300 VPWR.n206 VPWR.n198 0.120292
R3301 VPWR.n221 VPWR.n199 0.120292
R3302 VPWR.n216 VPWR.n199 0.120292
R3303 VPWR.n216 VPWR.n215 0.120292
R3304 VPWR.n215 VPWR.n214 0.120292
R3305 VPWR.n284 VPWR.n283 0.120292
R3306 VPWR.n285 VPWR.n284 0.120292
R3307 VPWR.n285 VPWR.n277 0.120292
R3308 VPWR.n300 VPWR.n278 0.120292
R3309 VPWR.n295 VPWR.n278 0.120292
R3310 VPWR.n295 VPWR.n294 0.120292
R3311 VPWR.n294 VPWR.n293 0.120292
R3312 VPWR.n124 VPWR.n123 0.120292
R3313 VPWR.n125 VPWR.n124 0.120292
R3314 VPWR.n125 VPWR.n117 0.120292
R3315 VPWR.n140 VPWR.n118 0.120292
R3316 VPWR.n135 VPWR.n118 0.120292
R3317 VPWR.n135 VPWR.n134 0.120292
R3318 VPWR.n134 VPWR.n133 0.120292
R3319 VPWR.n45 VPWR.n44 0.120292
R3320 VPWR.n46 VPWR.n45 0.120292
R3321 VPWR.n46 VPWR.n38 0.120292
R3322 VPWR.n61 VPWR.n39 0.120292
R3323 VPWR.n56 VPWR.n39 0.120292
R3324 VPWR.n56 VPWR.n55 0.120292
R3325 VPWR.n55 VPWR.n54 0.120292
R3326 VPWR.n422 VPWR.n421 0.120292
R3327 VPWR.n423 VPWR.n422 0.120292
R3328 VPWR.n423 VPWR.n415 0.120292
R3329 VPWR.n438 VPWR.n416 0.120292
R3330 VPWR.n433 VPWR.n416 0.120292
R3331 VPWR.n433 VPWR.n432 0.120292
R3332 VPWR.n432 VPWR.n431 0.120292
R3333 VPWR.n341 VPWR.n340 0.120292
R3334 VPWR.n342 VPWR.n341 0.120292
R3335 VPWR.n342 VPWR.n334 0.120292
R3336 VPWR.n357 VPWR.n335 0.120292
R3337 VPWR.n352 VPWR.n335 0.120292
R3338 VPWR.n352 VPWR.n351 0.120292
R3339 VPWR.n351 VPWR.n350 0.120292
R3340 VPWR.n584 VPWR.n583 0.120292
R3341 VPWR.n585 VPWR.n584 0.120292
R3342 VPWR.n585 VPWR.n577 0.120292
R3343 VPWR.n600 VPWR.n578 0.120292
R3344 VPWR.n595 VPWR.n578 0.120292
R3345 VPWR.n595 VPWR.n594 0.120292
R3346 VPWR.n594 VPWR.n593 0.120292
R3347 VPWR.n503 VPWR.n502 0.120292
R3348 VPWR.n504 VPWR.n503 0.120292
R3349 VPWR.n504 VPWR.n496 0.120292
R3350 VPWR.n519 VPWR.n497 0.120292
R3351 VPWR.n514 VPWR.n497 0.120292
R3352 VPWR.n514 VPWR.n513 0.120292
R3353 VPWR.n513 VPWR.n512 0.120292
R3354 VPWR.n222 VPWR.n221 0.115083
R3355 VPWR.n301 VPWR.n300 0.115083
R3356 VPWR.n141 VPWR.n140 0.115083
R3357 VPWR.n62 VPWR.n61 0.115083
R3358 VPWR.n439 VPWR.n438 0.115083
R3359 VPWR.n358 VPWR.n357 0.115083
R3360 VPWR.n601 VPWR.n600 0.115083
R3361 VPWR.n520 VPWR.n519 0.115083
R3362 VPWR.n414 VPWR 0.111772
R3363 VPWR VPWR.n560 0.109383
R3364 VPWR VPWR.n641 0.109383
R3365 VPWR.n196 VPWR.n195 0.0948367
R3366 VPWR.n275 VPWR.n274 0.0948367
R3367 VPWR.n115 VPWR.n114 0.0948367
R3368 VPWR.n36 VPWR.n35 0.0948367
R3369 VPWR.n477 VPWR.n476 0.0948367
R3370 VPWR.n396 VPWR.n395 0.0948367
R3371 VPWR.n639 VPWR.n638 0.0948367
R3372 VPWR.n558 VPWR.n557 0.0948367
R3373 VPWR VPWR.n398 0.0821625
R3374 VPWR VPWR.n479 0.0821625
R3375 VPWR.n196 VPWR.n180 0.0691538
R3376 VPWR.n275 VPWR.n259 0.0691538
R3377 VPWR.n115 VPWR.n99 0.0691538
R3378 VPWR.n36 VPWR.n20 0.0691538
R3379 VPWR.n477 VPWR.n461 0.0691538
R3380 VPWR.n396 VPWR.n380 0.0691538
R3381 VPWR.n639 VPWR.n623 0.0691538
R3382 VPWR.n558 VPWR.n542 0.0691538
R3383 VPWR.n197 VPWR.n196 0.0614341
R3384 VPWR.n276 VPWR.n275 0.0614341
R3385 VPWR.n116 VPWR.n115 0.0614341
R3386 VPWR.n37 VPWR.n36 0.0614341
R3387 VPWR.n478 VPWR.n477 0.0614341
R3388 VPWR.n397 VPWR.n396 0.0614341
R3389 VPWR.n640 VPWR.n639 0.0614341
R3390 VPWR.n559 VPWR.n558 0.0614341
R3391 VPWR.n158 VPWR 0.0613633
R3392 VPWR.n204 VPWR 0.0603958
R3393 VPWR.n283 VPWR 0.0603958
R3394 VPWR.n123 VPWR 0.0603958
R3395 VPWR.n44 VPWR 0.0603958
R3396 VPWR.n421 VPWR 0.0603958
R3397 VPWR.n340 VPWR 0.0603958
R3398 VPWR.n583 VPWR 0.0603958
R3399 VPWR.n502 VPWR 0.0603958
R3400 VPWR.n602 VPWR.n576 0.0565083
R3401 VPWR.n197 VPWR 0.0562442
R3402 VPWR.n276 VPWR 0.0562442
R3403 VPWR.n116 VPWR 0.0562442
R3404 VPWR.n37 VPWR 0.0562442
R3405 VPWR.n478 VPWR 0.0562442
R3406 VPWR.n397 VPWR 0.0562442
R3407 VPWR.n640 VPWR 0.0562442
R3408 VPWR.n559 VPWR 0.0562442
R3409 VPWR.n318 VPWR 0.0512194
R3410 VPWR.n229 VPWR 0.0459545
R3411 VPWR.n236 VPWR 0.0459545
R3412 VPWR.n308 VPWR 0.0459545
R3413 VPWR.n315 VPWR 0.0459545
R3414 VPWR.n69 VPWR 0.0459545
R3415 VPWR.n76 VPWR 0.0459545
R3416 VPWR.n148 VPWR 0.0459545
R3417 VPWR.n155 VPWR 0.0459545
R3418 VPWR.n405 VPWR 0.0459545
R3419 VPWR.n412 VPWR 0.0459545
R3420 VPWR.n325 VPWR 0.0459545
R3421 VPWR.n332 VPWR 0.0459545
R3422 VPWR.n567 VPWR 0.0459545
R3423 VPWR.n574 VPWR 0.0459545
R3424 VPWR.n487 VPWR 0.0459545
R3425 VPWR.n494 VPWR 0.0459545
R3426 VPWR.n440 VPWR.n414 0.0425062
R3427 VPWR.n229 VPWR 0.0338333
R3428 VPWR.n236 VPWR 0.0338333
R3429 VPWR.n308 VPWR 0.0338333
R3430 VPWR.n315 VPWR 0.0338333
R3431 VPWR.n69 VPWR 0.0338333
R3432 VPWR.n76 VPWR 0.0338333
R3433 VPWR.n148 VPWR 0.0338333
R3434 VPWR.n155 VPWR 0.0338333
R3435 VPWR.n405 VPWR 0.0338333
R3436 VPWR.n412 VPWR 0.0338333
R3437 VPWR.n325 VPWR 0.0338333
R3438 VPWR.n332 VPWR 0.0338333
R3439 VPWR.n567 VPWR 0.0338333
R3440 VPWR.n574 VPWR 0.0338333
R3441 VPWR.n487 VPWR 0.0338333
R3442 VPWR.n494 VPWR 0.0338333
R3443 VPWR.n214 VPWR 0.0226354
R3444 VPWR.n293 VPWR 0.0226354
R3445 VPWR.n133 VPWR 0.0226354
R3446 VPWR.n54 VPWR 0.0226354
R3447 VPWR.n431 VPWR 0.0226354
R3448 VPWR.n350 VPWR 0.0226354
R3449 VPWR.n593 VPWR 0.0226354
R3450 VPWR.n512 VPWR 0.0226354
R3451 VPWR VPWR.n642 0.006375
R3452 VPWR.n78 VPWR.n37 0.00599114
R3453 VPWR.n157 VPWR.n116 0.00599114
R3454 VPWR.n317 VPWR.n276 0.00599114
R3455 VPWR.n238 VPWR.n197 0.00599114
R3456 VPWR.n398 VPWR.n397 0.00599114
R3457 VPWR.n479 VPWR.n478 0.00599114
R3458 VPWR.n560 VPWR.n559 0.00599114
R3459 VPWR.n641 VPWR.n640 0.00599114
R3460 VPWR.n222 VPWR.n198 0.00570833
R3461 VPWR.n301 VPWR.n277 0.00570833
R3462 VPWR.n141 VPWR.n117 0.00570833
R3463 VPWR.n62 VPWR.n38 0.00570833
R3464 VPWR.n439 VPWR.n415 0.00570833
R3465 VPWR.n358 VPWR.n334 0.00570833
R3466 VPWR.n601 VPWR.n577 0.00570833
R3467 VPWR.n520 VPWR.n496 0.00570833
R3468 VPWR.n480 VPWR 0.00490625
R3469 VPWR.n238 VPWR.n159 0.00211964
R3470 VPWR VPWR.n317 0.00099705
R3471 VPWR VPWR.n157 0.000861799
R3472 VPWR.n318 VPWR 0.000831367
R3473 VPWR.n158 VPWR 0.000770504
R3474 VPWR.n157 VPWR.n78 0.000763741
R3475 VPWR.n317 VPWR.n238 0.000628489
R3476 ui_in[6].n2 ui_in[6].t1 212.081
R3477 ui_in[6].n1 ui_in[6].t4 212.081
R3478 ui_in[6].n6 ui_in[6].t6 212.081
R3479 ui_in[6].n0 ui_in[6].t7 212.081
R3480 ui_in[6].n11 ui_in[6].t5 212.081
R3481 ui_in[6].n17 ui_in[6].t0 212.081
R3482 ui_in[6].n12 ui_in[6].t2 212.081
R3483 ui_in[6].n13 ui_in[6].t18 212.081
R3484 ui_in[6] ui_in[6].n14 163.264
R3485 ui_in[6].n16 ui_in[6].n15 152
R3486 ui_in[6].n19 ui_in[6].n18 152
R3487 ui_in[6].n10 ui_in[6].n9 152
R3488 ui_in[6].n8 ui_in[6].n7 152
R3489 ui_in[6].n5 ui_in[6].n4 152
R3490 ui_in[6] ui_in[6].n3 152
R3491 ui_in[6].n2 ui_in[6].t12 139.78
R3492 ui_in[6].n1 ui_in[6].t14 139.78
R3493 ui_in[6].n6 ui_in[6].t16 139.78
R3494 ui_in[6].n0 ui_in[6].t17 139.78
R3495 ui_in[6].n11 ui_in[6].t15 139.78
R3496 ui_in[6].n17 ui_in[6].t11 139.78
R3497 ui_in[6].n12 ui_in[6].t13 139.78
R3498 ui_in[6].n13 ui_in[6].t9 139.78
R3499 ui_in[6].n24 ui_in[6].t19 120.23
R3500 ui_in[6].n24 ui_in[6].t3 120.228
R3501 ui_in[6].n21 ui_in[6].t8 118.061
R3502 ui_in[6].n21 ui_in[6].t10 118.058
R3503 ui_in[6].n3 ui_in[6].n2 30.6732
R3504 ui_in[6].n3 ui_in[6].n1 30.6732
R3505 ui_in[6].n5 ui_in[6].n1 30.6732
R3506 ui_in[6].n6 ui_in[6].n5 30.6732
R3507 ui_in[6].n7 ui_in[6].n6 30.6732
R3508 ui_in[6].n7 ui_in[6].n0 30.6732
R3509 ui_in[6].n10 ui_in[6].n0 30.6732
R3510 ui_in[6].n11 ui_in[6].n10 30.6732
R3511 ui_in[6].n18 ui_in[6].n11 30.6732
R3512 ui_in[6].n18 ui_in[6].n17 30.6732
R3513 ui_in[6].n17 ui_in[6].n16 30.6732
R3514 ui_in[6].n16 ui_in[6].n12 30.6732
R3515 ui_in[6].n14 ui_in[6].n12 30.6732
R3516 ui_in[6].n14 ui_in[6].n13 30.6732
R3517 ui_in[6].n4 ui_in[6] 21.5045
R3518 ui_in[6].n8 ui_in[6] 19.4565
R3519 ui_in[6].n9 ui_in[6] 17.4085
R3520 ui_in[6].n15 ui_in[6] 13.3125
R3521 ui_in[6].n20 ui_in[6].n19 13.0565
R3522 ui_in[6].n15 ui_in[6] 10.2405
R3523 ui_in[6].n19 ui_in[6] 8.1925
R3524 ui_in[6].n9 ui_in[6] 6.1445
R3525 ui_in[6] ui_in[6].n8 4.0965
R3526 ui_in[6].n23 ui_in[6].n20 3.2054
R3527 ui_in[6].n20 ui_in[6] 2.3045
R3528 ui_in[6].n4 ui_in[6] 2.0485
R3529 ui_in[6].n22 ui_in[6].n21 0.528909
R3530 ui_in[6].n25 ui_in[6].n24 0.506182
R3531 ui_in[6].n26 ui_in[6].n25 0.42675
R3532 ui_in[6].n26 ui_in[6].n23 0.342556
R3533 ui_in[6].n23 ui_in[6].n22 0.3415
R3534 ui_in[6].n25 ui_in[6] 0.170955
R3535 ui_in[6].n22 ui_in[6] 0.148227
R3536 ui_in[6] ui_in[6].n26 0.01225
R3537 ui_in[3].n2 ui_in[3].t17 212.081
R3538 ui_in[3].n1 ui_in[3].t15 212.081
R3539 ui_in[3].n6 ui_in[3].t16 212.081
R3540 ui_in[3].n0 ui_in[3].t12 212.081
R3541 ui_in[3].n11 ui_in[3].t8 212.081
R3542 ui_in[3].n17 ui_in[3].t9 212.081
R3543 ui_in[3].n12 ui_in[3].t11 212.081
R3544 ui_in[3].n13 ui_in[3].t13 212.081
R3545 ui_in[3] ui_in[3].n14 163.264
R3546 ui_in[3].n16 ui_in[3].n15 152
R3547 ui_in[3].n19 ui_in[3].n18 152
R3548 ui_in[3].n10 ui_in[3].n9 152
R3549 ui_in[3].n8 ui_in[3].n7 152
R3550 ui_in[3].n5 ui_in[3].n4 152
R3551 ui_in[3] ui_in[3].n3 152
R3552 ui_in[3].n2 ui_in[3].t7 139.78
R3553 ui_in[3].n1 ui_in[3].t5 139.78
R3554 ui_in[3].n6 ui_in[3].t6 139.78
R3555 ui_in[3].n0 ui_in[3].t2 139.78
R3556 ui_in[3].n11 ui_in[3].t18 139.78
R3557 ui_in[3].n17 ui_in[3].t19 139.78
R3558 ui_in[3].n12 ui_in[3].t1 139.78
R3559 ui_in[3].n13 ui_in[3].t3 139.78
R3560 ui_in[3].n24 ui_in[3].t0 120.23
R3561 ui_in[3].n24 ui_in[3].t10 120.228
R3562 ui_in[3].n21 ui_in[3].t14 118.061
R3563 ui_in[3].n21 ui_in[3].t4 118.058
R3564 ui_in[3].n3 ui_in[3].n2 30.6732
R3565 ui_in[3].n3 ui_in[3].n1 30.6732
R3566 ui_in[3].n5 ui_in[3].n1 30.6732
R3567 ui_in[3].n6 ui_in[3].n5 30.6732
R3568 ui_in[3].n7 ui_in[3].n6 30.6732
R3569 ui_in[3].n7 ui_in[3].n0 30.6732
R3570 ui_in[3].n10 ui_in[3].n0 30.6732
R3571 ui_in[3].n11 ui_in[3].n10 30.6732
R3572 ui_in[3].n18 ui_in[3].n11 30.6732
R3573 ui_in[3].n18 ui_in[3].n17 30.6732
R3574 ui_in[3].n17 ui_in[3].n16 30.6732
R3575 ui_in[3].n16 ui_in[3].n12 30.6732
R3576 ui_in[3].n14 ui_in[3].n12 30.6732
R3577 ui_in[3].n14 ui_in[3].n13 30.6732
R3578 ui_in[3].n4 ui_in[3] 21.5045
R3579 ui_in[3].n8 ui_in[3] 19.4565
R3580 ui_in[3].n9 ui_in[3] 17.4085
R3581 ui_in[3].n15 ui_in[3] 13.3125
R3582 ui_in[3].n20 ui_in[3].n19 13.0565
R3583 ui_in[3].n15 ui_in[3] 10.2405
R3584 ui_in[3].n19 ui_in[3] 8.1925
R3585 ui_in[3].n9 ui_in[3] 6.1445
R3586 ui_in[3] ui_in[3].n8 4.0965
R3587 ui_in[3].n23 ui_in[3].n20 3.2054
R3588 ui_in[3].n20 ui_in[3] 2.3045
R3589 ui_in[3].n4 ui_in[3] 2.0485
R3590 ui_in[3].n22 ui_in[3].n21 0.528909
R3591 ui_in[3].n25 ui_in[3].n24 0.506182
R3592 ui_in[3].n26 ui_in[3].n25 0.42675
R3593 ui_in[3].n26 ui_in[3].n23 0.342556
R3594 ui_in[3].n23 ui_in[3].n22 0.3415
R3595 ui_in[3].n25 ui_in[3] 0.170955
R3596 ui_in[3].n22 ui_in[3] 0.148227
R3597 ui_in[3] ui_in[3].n26 0.01225
R3598 distortionUnit_5.IN.n4 distortionUnit_5.IN.t4 223.565
R3599 distortionUnit_5.IN.n7 distortionUnit_5.IN.t5 223.565
R3600 distortionUnit_5.IN.n14 distortionUnit_5.IN.n12 199.941
R3601 distortionUnit_5.IN.n21 distortionUnit_5.IN.n20 199.941
R3602 distortionUnit_5.IN.n0 distortionUnit_5.IN.t14 118.769
R3603 distortionUnit_5.IN.n3 distortionUnit_5.IN.t12 118.621
R3604 distortionUnit_5.IN.n2 distortionUnit_5.IN.t16 118.005
R3605 distortionUnit_5.IN.n1 distortionUnit_5.IN.t15 118.005
R3606 distortionUnit_5.IN.n0 distortionUnit_5.IN.t13 118.005
R3607 distortionUnit_5.IN.n6 distortionUnit_5.IN.n5 90.2112
R3608 distortionUnit_5.IN.n22 distortionUnit_5.IN.t8 83.7234
R3609 distortionUnit_5.IN.n19 distortionUnit_5.IN.t9 83.7234
R3610 distortionUnit_5.IN.n13 distortionUnit_5.IN.t1 83.7234
R3611 distortionUnit_5.IN.n15 distortionUnit_5.IN.t0 83.7234
R3612 distortionUnit_5.IN.n6 distortionUnit_5.IN.n4 66.2405
R3613 distortionUnit_5.IN.n7 distortionUnit_5.IN.n6 63.2157
R3614 distortionUnit_5.IN.n12 distortionUnit_5.IN.t7 28.5655
R3615 distortionUnit_5.IN.n12 distortionUnit_5.IN.t6 28.5655
R3616 distortionUnit_5.IN.n20 distortionUnit_5.IN.t3 28.5655
R3617 distortionUnit_5.IN.n20 distortionUnit_5.IN.t2 28.5655
R3618 distortionUnit_5.IN.n5 distortionUnit_5.IN.t10 17.4005
R3619 distortionUnit_5.IN.n5 distortionUnit_5.IN.t11 17.4005
R3620 distortionUnit_5.IN.n8 distortionUnit_5.IN.n4 5.54823
R3621 distortionUnit_5.IN.n8 distortionUnit_5.IN.n7 5.18686
R3622 distortionUnit_5.IN.n10 distortionUnit_5.IN 4.9113
R3623 distortionUnit_5.IN.n9 distortionUnit_5.IN 4.4438
R3624 distortionUnit_5.IN distortionUnit_5.IN.n3 2.77717
R3625 distortionUnit_5.IN.n1 distortionUnit_5.IN.n0 2.66195
R3626 distortionUnit_5.IN.n3 distortionUnit_5.IN.n2 1.71868
R3627 distortionUnit_5.IN.n17 distortionUnit_5.IN.n16 1.15259
R3628 distortionUnit_5.IN.n18 distortionUnit_5.IN.n17 0.938152
R3629 distortionUnit_5.IN.n2 distortionUnit_5.IN.n1 0.764886
R3630 distortionUnit_5.IN.n13 distortionUnit_5.IN.n11 0.5005
R3631 distortionUnit_5.IN.n16 distortionUnit_5.IN.n15 0.5005
R3632 distortionUnit_5.IN.n19 distortionUnit_5.IN.n18 0.5005
R3633 distortionUnit_5.IN.n23 distortionUnit_5.IN.n22 0.5005
R3634 distortionUnit_5.IN.n9 distortionUnit_5.IN 0.490406
R3635 distortionUnit_5.IN.n21 distortionUnit_5.IN.n19 0.478385
R3636 distortionUnit_5.IN.n15 distortionUnit_5.IN.n14 0.478385
R3637 distortionUnit_5.IN.n14 distortionUnit_5.IN.n13 0.478385
R3638 distortionUnit_5.IN.n22 distortionUnit_5.IN.n21 0.478385
R3639 distortionUnit_5.IN.n16 distortionUnit_5.IN.n11 0.364136
R3640 distortionUnit_5.IN.n23 distortionUnit_5.IN.n18 0.364136
R3641 distortionUnit_5.IN.n11 distortionUnit_5.IN 0.244818
R3642 distortionUnit_5.IN distortionUnit_5.IN.n8 0.244818
R3643 distortionUnit_5.IN distortionUnit_5.IN.n23 0.244818
R3644 distortionUnit_5.IN distortionUnit_5.IN.n10 0.150313
R3645 distortionUnit_5.IN.n10 distortionUnit_5.IN 0.024
R3646 distortionUnit_5.IN.n17 distortionUnit_5.IN 0.0137188
R3647 distortionUnit_5.IN distortionUnit_5.IN.n9 0.0129412
R3648 ui_in[7].n2 ui_in[7].t5 212.081
R3649 ui_in[7].n1 ui_in[7].t9 212.081
R3650 ui_in[7].n6 ui_in[7].t3 212.081
R3651 ui_in[7].n0 ui_in[7].t4 212.081
R3652 ui_in[7].n11 ui_in[7].t8 212.081
R3653 ui_in[7].n17 ui_in[7].t2 212.081
R3654 ui_in[7].n12 ui_in[7].t6 212.081
R3655 ui_in[7].n13 ui_in[7].t1 212.081
R3656 ui_in[7] ui_in[7].n14 163.264
R3657 ui_in[7].n16 ui_in[7].n15 152
R3658 ui_in[7].n19 ui_in[7].n18 152
R3659 ui_in[7].n10 ui_in[7].n9 152
R3660 ui_in[7].n8 ui_in[7].n7 152
R3661 ui_in[7].n5 ui_in[7].n4 152
R3662 ui_in[7] ui_in[7].n3 152
R3663 ui_in[7].n2 ui_in[7].t15 139.78
R3664 ui_in[7].n1 ui_in[7].t18 139.78
R3665 ui_in[7].n6 ui_in[7].t13 139.78
R3666 ui_in[7].n0 ui_in[7].t14 139.78
R3667 ui_in[7].n11 ui_in[7].t17 139.78
R3668 ui_in[7].n17 ui_in[7].t12 139.78
R3669 ui_in[7].n12 ui_in[7].t16 139.78
R3670 ui_in[7].n13 ui_in[7].t11 139.78
R3671 ui_in[7].n24 ui_in[7].t19 120.23
R3672 ui_in[7].n24 ui_in[7].t0 120.228
R3673 ui_in[7].n21 ui_in[7].t7 118.061
R3674 ui_in[7].n21 ui_in[7].t10 118.058
R3675 ui_in[7].n3 ui_in[7].n2 30.6732
R3676 ui_in[7].n3 ui_in[7].n1 30.6732
R3677 ui_in[7].n5 ui_in[7].n1 30.6732
R3678 ui_in[7].n6 ui_in[7].n5 30.6732
R3679 ui_in[7].n7 ui_in[7].n6 30.6732
R3680 ui_in[7].n7 ui_in[7].n0 30.6732
R3681 ui_in[7].n10 ui_in[7].n0 30.6732
R3682 ui_in[7].n11 ui_in[7].n10 30.6732
R3683 ui_in[7].n18 ui_in[7].n11 30.6732
R3684 ui_in[7].n18 ui_in[7].n17 30.6732
R3685 ui_in[7].n17 ui_in[7].n16 30.6732
R3686 ui_in[7].n16 ui_in[7].n12 30.6732
R3687 ui_in[7].n14 ui_in[7].n12 30.6732
R3688 ui_in[7].n14 ui_in[7].n13 30.6732
R3689 ui_in[7].n4 ui_in[7] 21.5045
R3690 ui_in[7].n8 ui_in[7] 19.4565
R3691 ui_in[7].n9 ui_in[7] 17.4085
R3692 ui_in[7].n15 ui_in[7] 13.3125
R3693 ui_in[7].n20 ui_in[7].n19 13.0565
R3694 ui_in[7].n15 ui_in[7] 10.2405
R3695 ui_in[7].n19 ui_in[7] 8.1925
R3696 ui_in[7].n9 ui_in[7] 6.1445
R3697 ui_in[7] ui_in[7].n8 4.0965
R3698 ui_in[7].n23 ui_in[7].n20 3.2054
R3699 ui_in[7].n20 ui_in[7] 2.3045
R3700 ui_in[7].n4 ui_in[7] 2.0485
R3701 ui_in[7].n22 ui_in[7].n21 0.528909
R3702 ui_in[7].n25 ui_in[7].n24 0.506182
R3703 ui_in[7].n26 ui_in[7].n25 0.42675
R3704 ui_in[7].n26 ui_in[7].n23 0.342556
R3705 ui_in[7].n23 ui_in[7].n22 0.3415
R3706 ui_in[7].n25 ui_in[7] 0.170955
R3707 ui_in[7].n22 ui_in[7] 0.148227
R3708 ui_in[7] ui_in[7].n26 0.01225
R3709 ua[1].n9 ua[1].n7 199.941
R3710 ua[1].n3 ua[1].n1 199.941
R3711 ua[1].n8 ua[1].t0 83.7234
R3712 ua[1].n10 ua[1].t1 83.7234
R3713 ua[1].n2 ua[1].t6 83.7234
R3714 ua[1].n4 ua[1].t7 83.7234
R3715 ua[1].n7 ua[1].t4 28.5655
R3716 ua[1].n7 ua[1].t5 28.5655
R3717 ua[1].n1 ua[1].t3 28.5655
R3718 ua[1].n1 ua[1].t2 28.5655
R3719 ua[1].n13 ua[1] 4.9995
R3720 ua[1].n12 ua[1].n5 1.15259
R3721 ua[1].n12 ua[1].n11 0.938152
R3722 ua[1].n8 ua[1].n6 0.5005
R3723 ua[1].n11 ua[1].n10 0.5005
R3724 ua[1].n2 ua[1].n0 0.5005
R3725 ua[1].n5 ua[1].n4 0.5005
R3726 ua[1].n10 ua[1].n9 0.478385
R3727 ua[1].n9 ua[1].n8 0.478385
R3728 ua[1].n4 ua[1].n3 0.478385
R3729 ua[1].n3 ua[1].n2 0.478385
R3730 ua[1].n11 ua[1].n6 0.364136
R3731 ua[1].n5 ua[1].n0 0.364136
R3732 ua[1].n6 ua[1] 0.244818
R3733 ua[1].n0 ua[1] 0.244818
R3734 ua[1].n13 ua[1] 0.150313
R3735 ua[1] ua[1].n13 0.024
R3736 ua[1] ua[1].n12 0.0137188
R3737 ua[0].n4 ua[0].t0 223.565
R3738 ua[0].n7 ua[0].t1 223.565
R3739 ua[0].n0 ua[0].t4 118.769
R3740 ua[0].n3 ua[0].t7 118.621
R3741 ua[0].n2 ua[0].t5 118.005
R3742 ua[0].n1 ua[0].t6 118.005
R3743 ua[0].n0 ua[0].t8 118.005
R3744 ua[0].n6 ua[0].n5 90.2112
R3745 ua[0].n6 ua[0].n4 66.2405
R3746 ua[0].n7 ua[0].n6 63.2157
R3747 ua[0].n5 ua[0].t2 17.4005
R3748 ua[0].n5 ua[0].t3 17.4005
R3749 ua[0].n8 ua[0].n4 5.54823
R3750 ua[0].n8 ua[0].n7 5.18686
R3751 ua[0].n10 ua[0] 4.9402
R3752 ua[0].n9 ua[0] 4.4438
R3753 ua[0] ua[0].n10 3.53725
R3754 ua[0].n11 ua[0] 3.12125
R3755 ua[0] ua[0].n3 2.77717
R3756 ua[0].n1 ua[0].n0 2.66195
R3757 ua[0].n3 ua[0].n2 1.71868
R3758 ua[0].n2 ua[0].n1 0.764886
R3759 ua[0] ua[0].n8 0.244818
R3760 ua[0].n10 ua[0].n9 0.0729819
R3761 ua[0].n11 ua[0] 0.0480663
R3762 ua[0] ua[0].n11 0.0192548
R3763 ua[0].n9 ua[0] 0.013241
R3764 ui_in[2].n2 ui_in[2].t5 212.081
R3765 ui_in[2].n1 ui_in[2].t1 212.081
R3766 ui_in[2].n6 ui_in[2].t10 212.081
R3767 ui_in[2].n0 ui_in[2].t4 212.081
R3768 ui_in[2].n11 ui_in[2].t9 212.081
R3769 ui_in[2].n17 ui_in[2].t3 212.081
R3770 ui_in[2].n12 ui_in[2].t0 212.081
R3771 ui_in[2].n13 ui_in[2].t2 212.081
R3772 ui_in[2] ui_in[2].n14 163.264
R3773 ui_in[2].n16 ui_in[2].n15 152
R3774 ui_in[2].n19 ui_in[2].n18 152
R3775 ui_in[2].n10 ui_in[2].n9 152
R3776 ui_in[2].n8 ui_in[2].n7 152
R3777 ui_in[2].n5 ui_in[2].n4 152
R3778 ui_in[2] ui_in[2].n3 152
R3779 ui_in[2].n2 ui_in[2].t13 139.78
R3780 ui_in[2].n1 ui_in[2].t7 139.78
R3781 ui_in[2].n6 ui_in[2].t16 139.78
R3782 ui_in[2].n0 ui_in[2].t12 139.78
R3783 ui_in[2].n11 ui_in[2].t15 139.78
R3784 ui_in[2].n17 ui_in[2].t11 139.78
R3785 ui_in[2].n12 ui_in[2].t6 139.78
R3786 ui_in[2].n13 ui_in[2].t8 139.78
R3787 ui_in[2].n24 ui_in[2].t14 120.23
R3788 ui_in[2].n24 ui_in[2].t17 120.228
R3789 ui_in[2].n21 ui_in[2].t18 118.061
R3790 ui_in[2].n21 ui_in[2].t19 118.058
R3791 ui_in[2].n3 ui_in[2].n2 30.6732
R3792 ui_in[2].n3 ui_in[2].n1 30.6732
R3793 ui_in[2].n5 ui_in[2].n1 30.6732
R3794 ui_in[2].n6 ui_in[2].n5 30.6732
R3795 ui_in[2].n7 ui_in[2].n6 30.6732
R3796 ui_in[2].n7 ui_in[2].n0 30.6732
R3797 ui_in[2].n10 ui_in[2].n0 30.6732
R3798 ui_in[2].n11 ui_in[2].n10 30.6732
R3799 ui_in[2].n18 ui_in[2].n11 30.6732
R3800 ui_in[2].n18 ui_in[2].n17 30.6732
R3801 ui_in[2].n17 ui_in[2].n16 30.6732
R3802 ui_in[2].n16 ui_in[2].n12 30.6732
R3803 ui_in[2].n14 ui_in[2].n12 30.6732
R3804 ui_in[2].n14 ui_in[2].n13 30.6732
R3805 ui_in[2].n4 ui_in[2] 21.5045
R3806 ui_in[2].n8 ui_in[2] 19.4565
R3807 ui_in[2].n9 ui_in[2] 17.4085
R3808 ui_in[2].n15 ui_in[2] 13.3125
R3809 ui_in[2].n20 ui_in[2].n19 13.0565
R3810 ui_in[2].n15 ui_in[2] 10.2405
R3811 ui_in[2].n19 ui_in[2] 8.1925
R3812 ui_in[2].n9 ui_in[2] 6.1445
R3813 ui_in[2] ui_in[2].n8 4.0965
R3814 ui_in[2].n23 ui_in[2].n20 3.2054
R3815 ui_in[2].n20 ui_in[2] 2.3045
R3816 ui_in[2].n4 ui_in[2] 2.0485
R3817 ui_in[2].n22 ui_in[2].n21 0.528909
R3818 ui_in[2].n25 ui_in[2].n24 0.506182
R3819 ui_in[2].n26 ui_in[2].n25 0.42675
R3820 ui_in[2].n26 ui_in[2].n23 0.342556
R3821 ui_in[2].n23 ui_in[2].n22 0.3415
R3822 ui_in[2].n25 ui_in[2] 0.170955
R3823 ui_in[2].n22 ui_in[2] 0.148227
R3824 ui_in[2] ui_in[2].n26 0.01225
R3825 ui_in[5].n2 ui_in[5].t19 212.081
R3826 ui_in[5].n1 ui_in[5].t0 212.081
R3827 ui_in[5].n6 ui_in[5].t18 212.081
R3828 ui_in[5].n0 ui_in[5].t14 212.081
R3829 ui_in[5].n11 ui_in[5].t16 212.081
R3830 ui_in[5].n17 ui_in[5].t11 212.081
R3831 ui_in[5].n12 ui_in[5].t12 212.081
R3832 ui_in[5].n13 ui_in[5].t15 212.081
R3833 ui_in[5] ui_in[5].n14 163.264
R3834 ui_in[5].n16 ui_in[5].n15 152
R3835 ui_in[5].n19 ui_in[5].n18 152
R3836 ui_in[5].n10 ui_in[5].n9 152
R3837 ui_in[5].n8 ui_in[5].n7 152
R3838 ui_in[5].n5 ui_in[5].n4 152
R3839 ui_in[5] ui_in[5].n3 152
R3840 ui_in[5].n2 ui_in[5].t9 139.78
R3841 ui_in[5].n1 ui_in[5].t10 139.78
R3842 ui_in[5].n6 ui_in[5].t8 139.78
R3843 ui_in[5].n0 ui_in[5].t5 139.78
R3844 ui_in[5].n11 ui_in[5].t7 139.78
R3845 ui_in[5].n17 ui_in[5].t2 139.78
R3846 ui_in[5].n12 ui_in[5].t3 139.78
R3847 ui_in[5].n13 ui_in[5].t6 139.78
R3848 ui_in[5].n24 ui_in[5].t17 120.23
R3849 ui_in[5].n24 ui_in[5].t13 120.228
R3850 ui_in[5].n21 ui_in[5].t4 118.061
R3851 ui_in[5].n21 ui_in[5].t1 118.058
R3852 ui_in[5].n3 ui_in[5].n2 30.6732
R3853 ui_in[5].n3 ui_in[5].n1 30.6732
R3854 ui_in[5].n5 ui_in[5].n1 30.6732
R3855 ui_in[5].n6 ui_in[5].n5 30.6732
R3856 ui_in[5].n7 ui_in[5].n6 30.6732
R3857 ui_in[5].n7 ui_in[5].n0 30.6732
R3858 ui_in[5].n10 ui_in[5].n0 30.6732
R3859 ui_in[5].n11 ui_in[5].n10 30.6732
R3860 ui_in[5].n18 ui_in[5].n11 30.6732
R3861 ui_in[5].n18 ui_in[5].n17 30.6732
R3862 ui_in[5].n17 ui_in[5].n16 30.6732
R3863 ui_in[5].n16 ui_in[5].n12 30.6732
R3864 ui_in[5].n14 ui_in[5].n12 30.6732
R3865 ui_in[5].n14 ui_in[5].n13 30.6732
R3866 ui_in[5].n4 ui_in[5] 21.5045
R3867 ui_in[5].n8 ui_in[5] 19.4565
R3868 ui_in[5].n9 ui_in[5] 17.4085
R3869 ui_in[5].n15 ui_in[5] 13.3125
R3870 ui_in[5].n20 ui_in[5].n19 13.0565
R3871 ui_in[5].n15 ui_in[5] 10.2405
R3872 ui_in[5].n19 ui_in[5] 8.1925
R3873 ui_in[5].n9 ui_in[5] 6.1445
R3874 ui_in[5] ui_in[5].n8 4.0965
R3875 ui_in[5].n23 ui_in[5].n20 3.2054
R3876 ui_in[5].n20 ui_in[5] 2.3045
R3877 ui_in[5].n4 ui_in[5] 2.0485
R3878 ui_in[5].n22 ui_in[5].n21 0.528909
R3879 ui_in[5].n25 ui_in[5].n24 0.506182
R3880 ui_in[5].n26 ui_in[5].n25 0.42675
R3881 ui_in[5].n26 ui_in[5].n23 0.342556
R3882 ui_in[5].n23 ui_in[5].n22 0.3415
R3883 ui_in[5].n25 ui_in[5] 0.170955
R3884 ui_in[5].n22 ui_in[5] 0.148227
R3885 ui_in[5] ui_in[5].n26 0.01225
R3886 ui_in[1].n2 ui_in[1].t8 212.081
R3887 ui_in[1].n1 ui_in[1].t11 212.081
R3888 ui_in[1].n6 ui_in[1].t7 212.081
R3889 ui_in[1].n0 ui_in[1].t4 212.081
R3890 ui_in[1].n11 ui_in[1].t10 212.081
R3891 ui_in[1].n17 ui_in[1].t6 212.081
R3892 ui_in[1].n12 ui_in[1].t9 212.081
R3893 ui_in[1].n13 ui_in[1].t5 212.081
R3894 ui_in[1] ui_in[1].n14 163.264
R3895 ui_in[1].n16 ui_in[1].n15 152
R3896 ui_in[1].n19 ui_in[1].n18 152
R3897 ui_in[1].n10 ui_in[1].n9 152
R3898 ui_in[1].n8 ui_in[1].n7 152
R3899 ui_in[1].n5 ui_in[1].n4 152
R3900 ui_in[1] ui_in[1].n3 152
R3901 ui_in[1].n2 ui_in[1].t18 139.78
R3902 ui_in[1].n1 ui_in[1].t2 139.78
R3903 ui_in[1].n6 ui_in[1].t17 139.78
R3904 ui_in[1].n0 ui_in[1].t12 139.78
R3905 ui_in[1].n11 ui_in[1].t1 139.78
R3906 ui_in[1].n17 ui_in[1].t16 139.78
R3907 ui_in[1].n12 ui_in[1].t19 139.78
R3908 ui_in[1].n13 ui_in[1].t13 139.78
R3909 ui_in[1].n24 ui_in[1].t0 120.23
R3910 ui_in[1].n24 ui_in[1].t3 120.228
R3911 ui_in[1].n21 ui_in[1].t14 118.061
R3912 ui_in[1].n21 ui_in[1].t15 118.058
R3913 ui_in[1].n3 ui_in[1].n2 30.6732
R3914 ui_in[1].n3 ui_in[1].n1 30.6732
R3915 ui_in[1].n5 ui_in[1].n1 30.6732
R3916 ui_in[1].n6 ui_in[1].n5 30.6732
R3917 ui_in[1].n7 ui_in[1].n6 30.6732
R3918 ui_in[1].n7 ui_in[1].n0 30.6732
R3919 ui_in[1].n10 ui_in[1].n0 30.6732
R3920 ui_in[1].n11 ui_in[1].n10 30.6732
R3921 ui_in[1].n18 ui_in[1].n11 30.6732
R3922 ui_in[1].n18 ui_in[1].n17 30.6732
R3923 ui_in[1].n17 ui_in[1].n16 30.6732
R3924 ui_in[1].n16 ui_in[1].n12 30.6732
R3925 ui_in[1].n14 ui_in[1].n12 30.6732
R3926 ui_in[1].n14 ui_in[1].n13 30.6732
R3927 ui_in[1].n4 ui_in[1] 21.5045
R3928 ui_in[1].n8 ui_in[1] 19.4565
R3929 ui_in[1].n9 ui_in[1] 17.4085
R3930 ui_in[1].n15 ui_in[1] 13.3125
R3931 ui_in[1].n20 ui_in[1].n19 13.0565
R3932 ui_in[1].n15 ui_in[1] 10.2405
R3933 ui_in[1].n19 ui_in[1] 8.1925
R3934 ui_in[1].n9 ui_in[1] 6.1445
R3935 ui_in[1] ui_in[1].n8 4.0965
R3936 ui_in[1].n23 ui_in[1].n20 3.2054
R3937 ui_in[1].n20 ui_in[1] 2.3045
R3938 ui_in[1].n4 ui_in[1] 2.0485
R3939 ui_in[1].n22 ui_in[1].n21 0.528909
R3940 ui_in[1].n25 ui_in[1].n24 0.506182
R3941 ui_in[1].n26 ui_in[1].n25 0.42675
R3942 ui_in[1].n26 ui_in[1].n23 0.342556
R3943 ui_in[1].n23 ui_in[1].n22 0.3415
R3944 ui_in[1].n25 ui_in[1] 0.170955
R3945 ui_in[1].n22 ui_in[1] 0.148227
R3946 ui_in[1] ui_in[1].n26 0.01225
R3947 ui_in[0].n2 ui_in[0].t13 212.081
R3948 ui_in[0].n1 ui_in[0].t8 212.081
R3949 ui_in[0].n6 ui_in[0].t3 212.081
R3950 ui_in[0].n0 ui_in[0].t6 212.081
R3951 ui_in[0].n11 ui_in[0].t1 212.081
R3952 ui_in[0].n17 ui_in[0].t12 212.081
R3953 ui_in[0].n12 ui_in[0].t5 212.081
R3954 ui_in[0].n13 ui_in[0].t0 212.081
R3955 ui_in[0] ui_in[0].n14 163.264
R3956 ui_in[0].n16 ui_in[0].n15 152
R3957 ui_in[0].n19 ui_in[0].n18 152
R3958 ui_in[0].n10 ui_in[0].n9 152
R3959 ui_in[0].n8 ui_in[0].n7 152
R3960 ui_in[0].n5 ui_in[0].n4 152
R3961 ui_in[0] ui_in[0].n3 152
R3962 ui_in[0].n2 ui_in[0].t18 139.78
R3963 ui_in[0].n1 ui_in[0].t16 139.78
R3964 ui_in[0].n6 ui_in[0].t11 139.78
R3965 ui_in[0].n0 ui_in[0].t15 139.78
R3966 ui_in[0].n11 ui_in[0].t10 139.78
R3967 ui_in[0].n17 ui_in[0].t17 139.78
R3968 ui_in[0].n12 ui_in[0].t14 139.78
R3969 ui_in[0].n13 ui_in[0].t9 139.78
R3970 ui_in[0].n24 ui_in[0].t4 120.23
R3971 ui_in[0].n24 ui_in[0].t19 120.228
R3972 ui_in[0].n21 ui_in[0].t7 118.061
R3973 ui_in[0].n21 ui_in[0].t2 118.058
R3974 ui_in[0].n3 ui_in[0].n2 30.6732
R3975 ui_in[0].n3 ui_in[0].n1 30.6732
R3976 ui_in[0].n5 ui_in[0].n1 30.6732
R3977 ui_in[0].n6 ui_in[0].n5 30.6732
R3978 ui_in[0].n7 ui_in[0].n6 30.6732
R3979 ui_in[0].n7 ui_in[0].n0 30.6732
R3980 ui_in[0].n10 ui_in[0].n0 30.6732
R3981 ui_in[0].n11 ui_in[0].n10 30.6732
R3982 ui_in[0].n18 ui_in[0].n11 30.6732
R3983 ui_in[0].n18 ui_in[0].n17 30.6732
R3984 ui_in[0].n17 ui_in[0].n16 30.6732
R3985 ui_in[0].n16 ui_in[0].n12 30.6732
R3986 ui_in[0].n14 ui_in[0].n12 30.6732
R3987 ui_in[0].n14 ui_in[0].n13 30.6732
R3988 ui_in[0].n4 ui_in[0] 21.5045
R3989 ui_in[0].n8 ui_in[0] 19.4565
R3990 ui_in[0].n9 ui_in[0] 17.4085
R3991 ui_in[0].n15 ui_in[0] 13.3125
R3992 ui_in[0].n20 ui_in[0].n19 13.0565
R3993 ui_in[0].n15 ui_in[0] 10.2405
R3994 ui_in[0].n19 ui_in[0] 8.1925
R3995 ui_in[0].n9 ui_in[0] 6.1445
R3996 ui_in[0] ui_in[0].n8 4.0965
R3997 ui_in[0].n23 ui_in[0].n20 3.2054
R3998 ui_in[0].n20 ui_in[0] 2.3045
R3999 ui_in[0].n4 ui_in[0] 2.0485
R4000 ui_in[0].n22 ui_in[0].n21 0.528909
R4001 ui_in[0].n25 ui_in[0].n24 0.506182
R4002 ui_in[0].n26 ui_in[0].n25 0.42675
R4003 ui_in[0].n26 ui_in[0].n23 0.342556
R4004 ui_in[0].n23 ui_in[0].n22 0.3415
R4005 ui_in[0].n25 ui_in[0] 0.170955
R4006 ui_in[0].n22 ui_in[0] 0.148227
R4007 ui_in[0] ui_in[0].n26 0.01225
C0 distortionUnit_0.tgate_1.IN a_6908_16352# 0.001336f
C1 distortionUnit_5.IN distortionUnit_5.tgate_1.CTRLB 0.258603f
C2 a_7756_30557# distortionUnit_3.IN 3.11184f
C3 a_8010_16807# a_6908_16352# 1.5318f
C4 a_7876_23853# a_7032_23398# 0.27522f
C5 distortionUnit_5.tgate_1.IN a_8134_23853# 0.662032f
C6 ui_in[0] ui_in[7] 0.089842f
C7 distortionUnit_7.tgate_1.CTRLB distortionUnit_7.myOpamp_0.INn 9.97e-19
C8 distortionUnit_7.IN a_21192_16677# 0.763261f
C9 distortionUnit_7.tgate_1.CTRLB VPWR 4.29809f
C10 distortionUnit_5.IN distortionUnit_6.IN 1.38229f
C11 distortionUnit_7.sky130_fd_sc_hd__tap_2_0.VPB ui_in[7] 0.278876f
C12 distortionUnit_3.tgate_1.CTRLB ui_in[2] 2.30483f
C13 distortionUnit_3.IN a_6912_30102# 0.198383f
C14 distortionUnit_5.tgate_1.IN distortionUnit_5.myOpamp_0.INn 1.8069f
C15 distortionUnit_7.IN distortionUnit_7.myOpamp_0.INn 0.503808f
C16 ui_in[5] distortionUnit_6.sky130_fd_sc_hd__tap_2_0.VPB 0.278876f
C17 distortionUnit_2.IN distortionUnit_2.tgate_1.IN 0.820736f
C18 distortionUnit_2.IN distortionUnit_3.IN 1.3678f
C19 distortionUnit_0.myOpamp_0.INn distortionUnit_6.OUT 0.503808f
C20 VPWR distortionUnit_7.IN 12.891001f
C21 distortionUnit_5.tgate_1.IN ui_in[4] 0.795971f
C22 distortionUnit_2.IN ui_in[5] 0.238698f
C23 distortionUnit_1.sky130_fd_sc_hd__tap_2_0.VPB distortionUnit_3.IN 0.001709f
C24 distortionUnit_1.tgate_1.CTRLB distortionUnit_2.IN 1.62697f
C25 distortionUnit_2.IN ui_in[1] 1.59433f
C26 distortionUnit_3.tgate_1.IN distortionUnit_3.tgate_1.CTRLB 1.18065f
C27 ui_in[0] distortionUnit_1.myOpamp_0.INn 0.25444f
C28 distortionUnit_0.myOpamp_0.INn a_9638_15108# 0.007465f
C29 a_7968_36445# a_7710_36445# 1.57848f
C30 a_7756_30557# VPWR 4.6075f
C31 distortionUnit_1.sky130_fd_sc_hd__tap_2_0.VPB distortionUnit_1.tgate_1.CTRLB 0.175567f
C32 distortionUnit_4.IN a_20746_30481# 0.763261f
C33 ui_in[5] distortionUnit_6.OUT 1.93164f
C34 distortionUnit_2.IN ui_in[3] 0.284299f
C35 distortionUnit_1.myOpamp_0.INn a_7710_36445# 0.849481f
C36 distortionUnit_5.IN distortionUnit_4.tgate_1.CTRLB 1.6595f
C37 distortionUnit_7.tgate_1.CTRLB distortionUnit_7.IN 0.258603f
C38 a_20584_23723# VPWR 4.82533f
C39 VPWR a_6912_30102# 0.124672f
C40 a_7032_23398# VPWR 0.185809f
C41 VPWR distortionUnit_6.sky130_fd_sc_hd__tap_2_0.VPB 0.274328f
C42 distortionUnit_6.myOpamp_0.INn ui_in[5] 0.25444f
C43 distortionUnit_4.tgate_1.CTRLB distortionUnit_4.myOpamp_0.INn 9.97e-19
C44 distortionUnit_2.IN VPWR 15.030399f
C45 distortionUnit_1.sky130_fd_sc_hd__tap_2_0.VPB VPWR 0.274328f
C46 distortionUnit_3.IN ui_in[0] 0.067086f
C47 ui_in[5] ui_in[0] 0.087906f
C48 VPWR distortionUnit_6.OUT 13.9941f
C49 distortionUnit_2.tgate_1.CTRLB distortionUnit_2.myOpamp_0.INn 9.97e-19
C50 distortionUnit_4.IN distortionUnit_4.tgate_1.IN 0.820736f
C51 distortionUnit_1.tgate_1.CTRLB ui_in[0] 2.30483f
C52 distortionUnit_6.IN ui_in[7] 0.267407f
C53 distortionUnit_0.tgate_1.CTRLB ui_in[6] 2.30483f
C54 a_6866_35990# distortionUnit_1.tgate_1.IN 0.001336f
C55 ui_in[0] ui_in[1] 4.72532f
C56 distortionUnit_5.myOpamp_0.INn a_8134_23853# 1.23683f
C57 distortionUnit_4.IN distortionUnit_3.myOpamp_0.INn 0.005273f
C58 ui_in[6] ui_in[2] 0.085933f
C59 ui_in[5] distortionUnit_6.tgate_1.CTRLB 2.30483f
C60 distortionUnit_6.myOpamp_0.INn VPWR 1.38015f
C61 a_9642_28858# a_6912_30102# 6.06e-20
C62 ui_in[0] ui_in[3] 0.089682f
C63 ui_in[6] ui_in[4] 3.36528f
C64 distortionUnit_3.tgate_1.IN a_8014_30557# 0.662032f
C65 a_7756_30557# a_6912_30102# 0.27522f
C66 a_20746_30481# VPWR 0.156113f
C67 ui_in[2] ui_in[4] 1.79375f
C68 distortionUnit_5.myOpamp_0.INn ui_in[4] 0.25444f
C69 ui_in[0] VPWR 5.35341f
C70 a_20934_16677# a_21192_16677# 1.57848f
C71 a_19740_23268# VPWR 0.120584f
C72 distortionUnit_4.tgate_1.CTRLB distortionUnit_4.sky130_fd_sc_hd__tap_2_0.VPB 0.175567f
C73 distortionUnit_3.tgate_1.IN ui_in[2] 0.795971f
C74 distortionUnit_7.IN distortionUnit_6.OUT 1.3678f
C75 distortionUnit_3.IN distortionUnit_3.myOpamp_0.INn 0.503808f
C76 ui_in[5] a_22374_28782# 5e-19
C77 VPWR a_7710_36445# 4.55037f
C78 VPWR distortionUnit_7.sky130_fd_sc_hd__tap_2_0.VPB 0.274328f
C79 VPWR distortionUnit_6.tgate_1.CTRLB 4.49268f
C80 distortionUnit_5.IN distortionUnit_3.tgate_1.CTRLB 0.028918f
C81 a_20934_16677# distortionUnit_7.myOpamp_0.INn 0.849481f
C82 distortionUnit_5.tgate_1.IN distortionUnit_5.IN 0.820736f
C83 a_20782_36601# a_19680_36146# 1.5318f
C84 VPWR a_20934_16677# 4.53263f
C85 distortionUnit_4.tgate_1.IN ui_in[3] 0.795971f
C86 ua[0] a_6866_35990# 0.198383f
C87 distortionUnit_1.sky130_fd_sc_hd__tap_2_0.VPB distortionUnit_2.IN 4.57e-19
C88 distortionUnit_7.tgate_1.CTRLB distortionUnit_7.sky130_fd_sc_hd__tap_2_0.VPB 0.175567f
C89 VPWR distortionUnit_4.tgate_1.IN 6.29038f
C90 a_9596_34746# a_6866_35990# 6.06e-20
C91 distortionUnit_6.sky130_fd_sc_hd__tap_2_0.VPB distortionUnit_6.OUT 0.001873f
C92 VPWR distortionUnit_5.sky130_fd_sc_hd__tap_2_0.VPB 0.274328f
C93 a_20782_36601# a_20524_36601# 1.57848f
C94 VPWR distortionUnit_3.myOpamp_0.INn 0.698154f
C95 ui_in[5] distortionUnit_6.IN 1.32192f
C96 a_20584_23723# distortionUnit_6.myOpamp_0.INn 0.849481f
C97 distortionUnit_4.IN distortionUnit_4.tgate_1.CTRLB 0.258603f
C98 a_7752_16807# distortionUnit_0.tgate_1.IN 2.35765f
C99 distortionUnit_7.tgate_1.IN a_20090_16222# 0.001336f
C100 a_20934_16677# distortionUnit_7.IN 3.11184f
C101 a_7752_16807# a_8010_16807# 1.57848f
C102 a_19680_36146# a_22410_34902# 6.06e-20
C103 distortionUnit_5.tgate_1.CTRLB VPWR 4.58466f
C104 distortionUnit_6.tgate_1.IN a_20842_23723# 0.662032f
C105 a_20584_23723# a_19740_23268# 0.27522f
C106 a_7968_36445# a_6866_35990# 1.5318f
C107 distortionUnit_6.myOpamp_0.INn distortionUnit_6.OUT 0.260919f
C108 distortionUnit_2.IN ui_in[0] 1.89413f
C109 VPWR distortionUnit_6.IN 14.791201f
C110 distortionUnit_1.sky130_fd_sc_hd__tap_2_0.VPB ui_in[0] 0.278876f
C111 distortionUnit_1.myOpamp_0.INn a_6866_35990# 1.1307f
C112 distortionUnit_6.sky130_fd_sc_hd__tap_2_0.VPB distortionUnit_6.tgate_1.CTRLB 0.175567f
C113 a_9642_28858# distortionUnit_3.myOpamp_0.INn 0.007465f
C114 a_8134_23853# distortionUnit_5.IN 0.763261f
C115 a_20782_36601# distortionUnit_2.myOpamp_0.INn 1.23683f
C116 distortionUnit_5.IN ui_in[6] 0.232865f
C117 a_19680_36146# distortionUnit_2.tgate_1.IN 0.001336f
C118 distortionUnit_0.tgate_1.IN distortionUnit_0.myOpamp_0.INn 1.8069f
C119 a_19680_36146# distortionUnit_3.IN 5.62e-21
C120 a_7756_30557# distortionUnit_3.myOpamp_0.INn 0.849481f
C121 distortionUnit_4.tgate_1.CTRLB ui_in[3] 2.30483f
C122 distortionUnit_7.tgate_1.IN ua[1] 1.38344f
C123 a_19740_23268# distortionUnit_6.OUT 1.03e-19
C124 distortionUnit_5.IN ui_in[2] 0.044883f
C125 distortionUnit_5.myOpamp_0.INn a_9762_22154# 0.007465f
C126 a_22820_14978# a_20090_16222# 6.06e-20
C127 distortionUnit_5.myOpamp_0.INn distortionUnit_5.IN 0.503808f
C128 distortionUnit_0.myOpamp_0.INn a_8010_16807# 1.23683f
C129 distortionUnit_6.OUT distortionUnit_6.tgate_1.CTRLB 1.66142f
C130 VPWR distortionUnit_0.sky130_fd_sc_hd__tap_2_0.VPB 0.274328f
C131 distortionUnit_5.IN ui_in[4] 1.59742f
C132 distortionUnit_6.myOpamp_0.INn a_19740_23268# 1.1307f
C133 VPWR distortionUnit_4.tgate_1.CTRLB 4.30804f
C134 distortionUnit_3.myOpamp_0.INn a_6912_30102# 1.1307f
C135 a_20524_36601# distortionUnit_2.tgate_1.IN 2.35765f
C136 distortionUnit_3.IN a_6866_35990# 6.34e-19
C137 distortionUnit_6.myOpamp_0.INn distortionUnit_6.tgate_1.CTRLB 9.97e-19
C138 distortionUnit_4.IN distortionUnit_3.tgate_1.CTRLB 1.62697f
C139 a_19680_36146# VPWR 0.138823f
C140 distortionUnit_5.sky130_fd_sc_hd__tap_2_0.VPB distortionUnit_6.OUT 0.001173f
C141 a_22410_34902# distortionUnit_2.myOpamp_0.INn 0.007465f
C142 ua[0] ua[1] 0.45455f
C143 a_7876_23853# distortionUnit_5.tgate_1.IN 2.35765f
C144 a_20584_23723# distortionUnit_6.IN 3.11184f
C145 distortionUnit_0.tgate_1.IN VPWR 6.9119f
C146 distortionUnit_7.IN distortionUnit_0.sky130_fd_sc_hd__tap_2_0.VPB 4.57e-19
C147 VPWR a_20524_36601# 4.64125f
C148 a_19644_30026# a_20488_30481# 0.27522f
C149 a_20746_30481# distortionUnit_4.tgate_1.IN 0.662032f
C150 distortionUnit_3.IN distortionUnit_3.tgate_1.CTRLB 0.258603f
C151 VPWR a_6866_35990# 0.100029f
C152 distortionUnit_5.tgate_1.CTRLB distortionUnit_6.OUT 0.028102f
C153 VPWR a_8010_16807# 0.156762f
C154 ui_in[6] ui_in[7] 7.30655f
C155 distortionUnit_2.tgate_1.IN distortionUnit_2.myOpamp_0.INn 1.8069f
C156 distortionUnit_3.IN distortionUnit_2.myOpamp_0.INn 0.23705f
C157 ui_in[7] ua[1] 1.87785f
C158 ui_in[2] ui_in[7] 0.086999f
C159 distortionUnit_6.IN distortionUnit_6.OUT 1.3678f
C160 ui_in[1] distortionUnit_2.myOpamp_0.INn 0.25444f
C161 ui_in[7] ui_in[4] 0.089626f
C162 distortionUnit_3.tgate_1.CTRLB distortionUnit_3.sky130_fd_sc_hd__tap_2_0.VPB 0.175567f
C163 distortionUnit_2.myOpamp_0.INn ui_in[3] 0.058805f
C164 distortionUnit_0.tgate_1.IN distortionUnit_7.IN 1.38344f
C165 distortionUnit_5.IN a_19644_30026# 5.62e-21
C166 distortionUnit_6.myOpamp_0.INn distortionUnit_6.IN 0.503808f
C167 distortionUnit_3.tgate_1.CTRLB VPWR 4.37242f
C168 distortionUnit_5.tgate_1.IN VPWR 7.473f
C169 a_20488_30481# distortionUnit_4.myOpamp_0.INn 0.849481f
C170 a_19644_30026# distortionUnit_4.myOpamp_0.INn 1.1307f
C171 VPWR distortionUnit_2.myOpamp_0.INn 0.867237f
C172 a_7752_16807# a_6908_16352# 0.27522f
C173 distortionUnit_4.IN ui_in[6] 0.244964f
C174 a_19680_36146# distortionUnit_2.IN 0.198383f
C175 a_21192_16677# a_20090_16222# 1.5318f
C176 a_19740_23268# distortionUnit_6.IN 0.198383f
C177 distortionUnit_4.IN ui_in[2] 1.89891f
C178 a_7876_23853# a_8134_23853# 1.57848f
C179 ui_in[6] distortionUnit_0.myOpamp_0.INn 0.25444f
C180 distortionUnit_0.tgate_1.CTRLB distortionUnit_0.myOpamp_0.INn 9.97e-19
C181 distortionUnit_6.IN distortionUnit_6.tgate_1.CTRLB 0.258603f
C182 distortionUnit_4.IN ui_in[4] 0.261488f
C183 distortionUnit_7.myOpamp_0.INn a_20090_16222# 1.1307f
C184 distortionUnit_5.IN distortionUnit_4.myOpamp_0.INn 0.236699f
C185 VPWR a_20090_16222# 0.100029f
C186 distortionUnit_3.IN a_8014_30557# 0.763261f
C187 a_7876_23853# distortionUnit_5.myOpamp_0.INn 0.849481f
C188 distortionUnit_3.tgate_1.IN distortionUnit_4.IN 1.38344f
C189 distortionUnit_3.IN ui_in[6] 0.234443f
C190 distortionUnit_2.IN a_20524_36601# 3.11184f
C191 ui_in[5] ui_in[6] 3.7149f
C192 distortionUnit_5.tgate_1.CTRLB distortionUnit_5.sky130_fd_sc_hd__tap_2_0.VPB 0.175567f
C193 distortionUnit_0.tgate_1.IN distortionUnit_6.OUT 0.820736f
C194 distortionUnit_3.IN ui_in[2] 1.74342f
C195 ui_in[6] ui_in[1] 0.17014f
C196 ui_in[5] ui_in[2] 0.086037f
C197 ua[0] distortionUnit_1.tgate_1.IN 0.820736f
C198 distortionUnit_0.myOpamp_0.INn a_6908_16352# 1.1307f
C199 distortionUnit_1.tgate_1.CTRLB ui_in[2] 0.005458f
C200 distortionUnit_5.sky130_fd_sc_hd__tap_2_0.VPB distortionUnit_6.IN 4.57e-19
C201 distortionUnit_3.IN ui_in[4] 0.234366f
C202 ui_in[1] ui_in[2] 4.51989f
C203 a_8010_16807# distortionUnit_6.OUT 0.763261f
C204 ui_in[6] ui_in[3] 0.166581f
C205 ui_in[5] ui_in[4] 3.90346f
C206 distortionUnit_3.tgate_1.IN distortionUnit_3.IN 0.820736f
C207 ui_in[2] ui_in[3] 3.92737f
C208 ui_in[1] ui_in[4] 0.174472f
C209 distortionUnit_5.tgate_1.IN a_7032_23398# 0.001336f
C210 VPWR a_8014_30557# 0.161318f
C211 a_8134_23853# VPWR 0.193581f
C212 distortionUnit_7.IN a_20090_16222# 0.198383f
C213 ui_in[2] distortionUnit_3.sky130_fd_sc_hd__tap_2_0.VPB 0.278876f
C214 ui_in[6] VPWR 5.42895f
C215 distortionUnit_7.myOpamp_0.INn ua[1] 0.005273f
C216 distortionUnit_0.tgate_1.CTRLB VPWR 4.4067f
C217 ui_in[3] ui_in[4] 3.73034f
C218 distortionUnit_5.tgate_1.CTRLB distortionUnit_6.IN 1.62697f
C219 VPWR ua[1] 3.53963f
C220 distortionUnit_6.tgate_1.IN ui_in[5] 0.795971f
C221 distortionUnit_4.tgate_1.CTRLB distortionUnit_4.tgate_1.IN 1.18065f
C222 distortionUnit_2.IN distortionUnit_2.myOpamp_0.INn 0.503808f
C223 VPWR ui_in[2] 5.62877f
C224 distortionUnit_5.myOpamp_0.INn VPWR 1.83805f
C225 distortionUnit_5.IN distortionUnit_4.sky130_fd_sc_hd__tap_2_0.VPB 0.001804f
C226 distortionUnit_5.IN ui_in[7] 0.238801f
C227 distortionUnit_7.tgate_1.IN ui_in[7] 0.795971f
C228 VPWR ui_in[4] 5.66871f
C229 distortionUnit_4.IN a_20488_30481# 3.11184f
C230 a_6866_35990# a_7710_36445# 0.27522f
C231 a_7968_36445# distortionUnit_1.tgate_1.IN 0.662032f
C232 distortionUnit_3.tgate_1.IN VPWR 6.64767f
C233 distortionUnit_2.tgate_1.CTRLB distortionUnit_2.tgate_1.IN 1.18065f
C234 distortionUnit_7.tgate_1.CTRLB ua[1] 1.62697f
C235 distortionUnit_3.IN distortionUnit_2.tgate_1.CTRLB 1.65953f
C236 distortionUnit_4.IN a_19644_30026# 0.198383f
C237 VPWR a_6908_16352# 0.100029f
C238 distortionUnit_1.myOpamp_0.INn distortionUnit_1.tgate_1.IN 1.8069f
C239 ui_in[6] distortionUnit_7.IN 1.90243f
C240 distortionUnit_6.tgate_1.IN VPWR 7.26402f
C241 ui_in[1] distortionUnit_2.tgate_1.CTRLB 2.30483f
C242 distortionUnit_0.tgate_1.CTRLB distortionUnit_7.IN 1.62697f
C243 distortionUnit_7.IN ua[1] 1.3678f
C244 a_7756_30557# a_8014_30557# 1.57848f
C245 distortionUnit_2.sky130_fd_sc_hd__tap_2_0.VPB distortionUnit_2.tgate_1.CTRLB 0.175567f
C246 distortionUnit_4.IN distortionUnit_5.IN 1.3678f
C247 a_20842_23723# VPWR 0.164659f
C248 a_8134_23853# a_7032_23398# 1.5318f
C249 a_8014_30557# a_6912_30102# 1.5318f
C250 VPWR distortionUnit_2.tgate_1.CTRLB 4.40906f
C251 distortionUnit_4.IN distortionUnit_4.myOpamp_0.INn 0.503808f
C252 a_7876_23853# distortionUnit_5.IN 3.11184f
C253 ua[0] a_7968_36445# 0.763261f
C254 distortionUnit_2.IN ui_in[6] 0.234969f
C255 a_7756_30557# distortionUnit_3.tgate_1.IN 2.35765f
C256 distortionUnit_5.myOpamp_0.INn a_7032_23398# 1.1307f
C257 distortionUnit_1.tgate_1.CTRLB distortionUnit_1.tgate_1.IN 1.18065f
C258 distortionUnit_5.IN distortionUnit_3.IN 0.185605f
C259 distortionUnit_2.IN ui_in[2] 0.262185f
C260 ua[0] distortionUnit_1.myOpamp_0.INn 0.503808f
C261 distortionUnit_5.IN ui_in[5] 0.337455f
C262 VPWR a_20488_30481# 4.57345f
C263 ui_in[6] distortionUnit_6.OUT 1.58548f
C264 distortionUnit_2.IN ui_in[4] 0.236324f
C265 distortionUnit_0.tgate_1.CTRLB distortionUnit_6.OUT 0.258603f
C266 distortionUnit_3.tgate_1.IN a_6912_30102# 0.001336f
C267 distortionUnit_3.tgate_1.CTRLB distortionUnit_3.myOpamp_0.INn 9.97e-19
C268 a_19644_30026# VPWR 0.101675f
C269 a_9596_34746# distortionUnit_1.myOpamp_0.INn 0.007465f
C270 ui_in[5] distortionUnit_4.myOpamp_0.INn 0.03372f
C271 a_20934_16677# a_20090_16222# 0.27522f
C272 distortionUnit_7.tgate_1.IN a_21192_16677# 0.662032f
C273 distortionUnit_5.IN ui_in[3] 1.92809f
C274 distortionUnit_5.myOpamp_0.INn distortionUnit_6.OUT 0.182465f
C275 a_20584_23723# distortionUnit_6.tgate_1.IN 2.35765f
C276 distortionUnit_5.IN distortionUnit_3.sky130_fd_sc_hd__tap_2_0.VPB 0.001206f
C277 distortionUnit_6.OUT ui_in[4] 0.043613f
C278 VPWR distortionUnit_1.tgate_1.IN 5.98641f
C279 distortionUnit_5.tgate_1.IN distortionUnit_5.tgate_1.CTRLB 1.18065f
C280 distortionUnit_7.tgate_1.IN distortionUnit_7.myOpamp_0.INn 1.8069f
C281 distortionUnit_4.myOpamp_0.INn ui_in[3] 0.25444f
C282 distortionUnit_5.IN VPWR 15.008401f
C283 VPWR distortionUnit_7.tgate_1.IN 6.25187f
C284 a_20584_23723# a_20842_23723# 1.57848f
C285 distortionUnit_4.IN ui_in[7] 0.253945f
C286 a_6908_16352# distortionUnit_6.OUT 0.198383f
C287 ui_in[6] ui_in[0] 0.088028f
C288 distortionUnit_5.tgate_1.IN distortionUnit_6.IN 1.38344f
C289 distortionUnit_1.tgate_1.CTRLB ua[0] 0.258603f
C290 VPWR distortionUnit_4.myOpamp_0.INn 0.578814f
C291 distortionUnit_6.tgate_1.IN distortionUnit_6.OUT 1.38344f
C292 ui_in[0] ui_in[2] 1.02988f
C293 distortionUnit_1.myOpamp_0.INn a_7968_36445# 1.23683f
C294 a_6908_16352# a_9638_15108# 6.06e-20
C295 distortionUnit_3.IN a_9596_34746# 0.023593f
C296 distortionUnit_2.IN distortionUnit_2.tgate_1.CTRLB 0.258603f
C297 distortionUnit_7.sky130_fd_sc_hd__tap_2_0.VPB ua[1] 4.57e-19
C298 ui_in[0] ui_in[4] 0.089269f
C299 a_19680_36146# a_20524_36601# 0.27522f
C300 a_7752_16807# distortionUnit_0.myOpamp_0.INn 0.849481f
C301 a_20782_36601# distortionUnit_2.tgate_1.IN 0.662032f
C302 distortionUnit_7.tgate_1.CTRLB distortionUnit_7.tgate_1.IN 1.18065f
C303 distortionUnit_6.tgate_1.IN distortionUnit_6.myOpamp_0.INn 1.8069f
C304 distortionUnit_3.IN ui_in[7] 0.240454f
C305 ui_in[5] ui_in[7] 2.54379f
C306 distortionUnit_5.IN a_9642_28858# 0.011741f
C307 ua[0] VPWR 20.3921f
C308 distortionUnit_7.tgate_1.IN distortionUnit_7.IN 0.820736f
C309 distortionUnit_0.tgate_1.IN a_8010_16807# 0.662032f
C310 ui_in[1] ui_in[7] 0.18869f
C311 distortionUnit_6.myOpamp_0.INn a_20842_23723# 1.23683f
C312 a_22820_14978# distortionUnit_7.myOpamp_0.INn 0.007465f
C313 distortionUnit_3.myOpamp_0.INn a_8014_30557# 1.23683f
C314 distortionUnit_6.tgate_1.IN a_19740_23268# 0.001336f
C315 distortionUnit_4.sky130_fd_sc_hd__tap_2_0.VPB ui_in[3] 0.278876f
C316 ui_in[7] ui_in[3] 0.184684f
C317 ui_in[2] distortionUnit_3.myOpamp_0.INn 0.25444f
C318 distortionUnit_6.tgate_1.IN distortionUnit_6.tgate_1.CTRLB 1.18065f
C319 a_20782_36601# VPWR 0.164599f
C320 distortionUnit_3.IN distortionUnit_1.myOpamp_0.INn 0.396323f
C321 distortionUnit_7.myOpamp_0.INn ui_in[7] 0.25444f
C322 a_7032_23398# a_9762_22154# 6.06e-20
C323 distortionUnit_5.sky130_fd_sc_hd__tap_2_0.VPB ui_in[4] 0.278876f
C324 distortionUnit_2.IN distortionUnit_1.tgate_1.IN 1.38344f
C325 a_7032_23398# distortionUnit_5.IN 0.198383f
C326 a_20842_23723# a_19740_23268# 1.5318f
C327 VPWR distortionUnit_4.sky130_fd_sc_hd__tap_2_0.VPB 0.274328f
C328 a_19680_36146# distortionUnit_2.myOpamp_0.INn 1.1307f
C329 VPWR ui_in[7] 5.46148f
C330 distortionUnit_1.tgate_1.CTRLB distortionUnit_1.myOpamp_0.INn 9.97e-19
C331 distortionUnit_4.IN distortionUnit_3.IN 1.61854f
C332 a_22410_34902# distortionUnit_3.IN 0.014606f
C333 distortionUnit_4.IN ui_in[5] 0.291464f
C334 distortionUnit_3.tgate_1.IN distortionUnit_3.myOpamp_0.INn 1.8069f
C335 a_7752_16807# VPWR 4.63532f
C336 a_22470_22024# distortionUnit_6.OUT 0.016146f
C337 distortionUnit_5.myOpamp_0.INn distortionUnit_5.tgate_1.CTRLB 9.97e-19
C338 ui_in[6] distortionUnit_6.IN 0.255482f
C339 a_20746_30481# a_20488_30481# 1.57848f
C340 distortionUnit_5.tgate_1.CTRLB ui_in[4] 2.30483f
C341 a_9762_22154# distortionUnit_6.OUT 0.011183f
C342 VPWR a_7968_36445# 0.150636f
C343 distortionUnit_6.myOpamp_0.INn a_22470_22024# 0.007465f
C344 distortionUnit_7.tgate_1.CTRLB ui_in[7] 2.30483f
C345 distortionUnit_4.IN ui_in[3] 1.31839f
C346 distortionUnit_5.myOpamp_0.INn distortionUnit_6.IN 0.005273f
C347 a_20524_36601# distortionUnit_2.myOpamp_0.INn 0.849481f
C348 a_22410_34902# ui_in[3] 0.001393f
C349 a_20746_30481# a_19644_30026# 1.5318f
C350 VPWR distortionUnit_1.myOpamp_0.INn 0.537507f
C351 distortionUnit_4.IN distortionUnit_3.sky130_fd_sc_hd__tap_2_0.VPB 4.57e-19
C352 distortionUnit_3.IN distortionUnit_2.tgate_1.IN 1.38344f
C353 distortionUnit_6.IN ui_in[4] 1.90075f
C354 distortionUnit_3.IN ui_in[5] 0.233538f
C355 distortionUnit_7.IN ui_in[7] 1.33097f
C356 distortionUnit_1.tgate_1.CTRLB distortionUnit_3.IN 0.043142f
C357 distortionUnit_4.IN VPWR 15.4213f
C358 ui_in[1] distortionUnit_2.tgate_1.IN 0.795971f
C359 ui_in[6] distortionUnit_0.sky130_fd_sc_hd__tap_2_0.VPB 0.278876f
C360 distortionUnit_3.IN ui_in[1] 1.92857f
C361 distortionUnit_2.IN ua[0] 1.3678f
C362 distortionUnit_0.tgate_1.CTRLB distortionUnit_0.sky130_fd_sc_hd__tap_2_0.VPB 0.175567f
C363 ui_in[5] ui_in[1] 0.172407f
C364 a_19740_23268# a_22470_22024# 6.06e-20
C365 ui_in[0] distortionUnit_1.tgate_1.IN 0.795971f
C366 distortionUnit_0.myOpamp_0.INn VPWR 0.878609f
C367 distortionUnit_2.sky130_fd_sc_hd__tap_2_0.VPB distortionUnit_3.IN 0.001804f
C368 distortionUnit_3.IN ui_in[3] 1.11357f
C369 distortionUnit_6.tgate_1.IN distortionUnit_6.IN 0.820736f
C370 ui_in[5] ui_in[3] 2.18372f
C371 a_7876_23853# VPWR 5.38803f
C372 a_7710_36445# distortionUnit_1.tgate_1.IN 2.35765f
C373 a_20488_30481# distortionUnit_4.tgate_1.IN 2.35765f
C374 a_20746_30481# distortionUnit_4.myOpamp_0.INn 1.23683f
C375 distortionUnit_2.sky130_fd_sc_hd__tap_2_0.VPB ui_in[1] 0.278876f
C376 ui_in[1] ui_in[3] 1.03886f
C377 a_19644_30026# distortionUnit_4.tgate_1.IN 0.001336f
C378 VPWR distortionUnit_2.tgate_1.IN 6.88843f
C379 a_20782_36601# distortionUnit_2.IN 0.763261f
C380 distortionUnit_3.IN VPWR 14.905f
C381 a_20842_23723# distortionUnit_6.IN 0.763261f
C382 ui_in[5] VPWR 5.68023f
C383 distortionUnit_2.IN ui_in[7] 0.24347f
C384 a_19644_30026# a_22374_28782# 6.06e-20
C385 a_20934_16677# distortionUnit_7.tgate_1.IN 2.35765f
C386 distortionUnit_1.tgate_1.CTRLB VPWR 4.27547f
C387 VPWR ui_in[1] 5.30897f
C388 ui_in[6] distortionUnit_0.tgate_1.IN 0.795971f
C389 distortionUnit_0.tgate_1.CTRLB distortionUnit_0.tgate_1.IN 1.18065f
C390 distortionUnit_7.myOpamp_0.INn a_21192_16677# 1.23683f
C391 VPWR a_21192_16677# 0.148886f
C392 distortionUnit_2.sky130_fd_sc_hd__tap_2_0.VPB VPWR 0.274328f
C393 VPWR ui_in[3] 5.65932f
C394 distortionUnit_5.IN distortionUnit_4.tgate_1.IN 1.38344f
C395 distortionUnit_6.OUT ui_in[7] 0.317052f
C396 distortionUnit_0.myOpamp_0.INn distortionUnit_7.IN 0.005273f
C397 ui_in[0] ua[0] 1.30899f
C398 VPWR distortionUnit_3.sky130_fd_sc_hd__tap_2_0.VPB 0.274328f
C399 distortionUnit_5.IN a_22374_28782# 0.014536f
C400 distortionUnit_5.IN distortionUnit_3.myOpamp_0.INn 0.190753f
C401 a_7752_16807# distortionUnit_6.OUT 3.11184f
C402 VPWR distortionUnit_7.myOpamp_0.INn 0.534285f
C403 distortionUnit_4.tgate_1.IN distortionUnit_4.myOpamp_0.INn 1.8069f
C404 ua[0] a_7710_36445# 3.11184f
C405 distortionUnit_2.IN distortionUnit_1.myOpamp_0.INn 0.005273f
C406 distortionUnit_6.myOpamp_0.INn ui_in[7] 0.030058f
C407 a_22374_28782# distortionUnit_4.myOpamp_0.INn 0.007465f
C408 ua[1] VGND 20.273489f
C409 ui_in[7] VGND 30.446981f
C410 ui_in[6] VGND 28.304464f
C411 ui_in[5] VGND 28.04565f
C412 ui_in[4] VGND 24.38021f
C413 ui_in[3] VGND 24.552017f
C414 ui_in[2] VGND 21.405964f
C415 ui_in[1] VGND 21.530247f
C416 ua[0] VGND 60.84894f
C417 ui_in[0] VGND 20.35954f
C418 VPWR VGND -0.241886p
C419 distortionUnit_7.tgate_1.CTRLB VGND 4.90769f
C420 a_22820_14978# VGND 0.672562f
C421 a_20090_16222# VGND 5.77883f
C422 a_21192_16677# VGND 1.79918f
C423 distortionUnit_7.myOpamp_0.INn VGND 8.781199f
C424 distortionUnit_7.tgate_1.IN VGND 2.92383f
C425 a_20934_16677# VGND 4.02935f
C426 distortionUnit_0.tgate_1.CTRLB VGND 4.92215f
C427 a_9638_15108# VGND 0.673165f
C428 a_6908_16352# VGND 5.7588f
C429 a_8010_16807# VGND 1.78029f
C430 distortionUnit_0.myOpamp_0.INn VGND 8.510679f
C431 distortionUnit_0.tgate_1.IN VGND 2.6941f
C432 a_7752_16807# VGND 3.58914f
C433 distortionUnit_7.IN VGND 14.596201f
C434 distortionUnit_6.tgate_1.CTRLB VGND 4.86682f
C435 a_22470_22024# VGND 0.673612f
C436 a_19740_23268# VGND 5.71223f
C437 a_20842_23723# VGND 1.74561f
C438 distortionUnit_6.myOpamp_0.INn VGND 8.04186f
C439 distortionUnit_6.tgate_1.IN VGND 2.59761f
C440 a_20584_23723# VGND 3.11162f
C441 distortionUnit_5.tgate_1.CTRLB VGND 4.79446f
C442 a_9762_22154# VGND 0.680066f
C443 a_7032_23398# VGND 5.62738f
C444 a_8134_23853# VGND 1.69448f
C445 distortionUnit_5.myOpamp_0.INn VGND 8.043759f
C446 distortionUnit_5.tgate_1.IN VGND 2.55687f
C447 a_7876_23853# VGND 2.82463f
C448 distortionUnit_6.OUT VGND 30.295801f
C449 distortionUnit_6.IN VGND 13.4661f
C450 distortionUnit_4.tgate_1.CTRLB VGND 4.89096f
C451 a_22374_28782# VGND 0.673472f
C452 a_19644_30026# VGND 5.73689f
C453 a_20746_30481# VGND 1.75741f
C454 distortionUnit_4.myOpamp_0.INn VGND 8.11164f
C455 distortionUnit_4.tgate_1.IN VGND 2.68792f
C456 a_20488_30481# VGND 3.28069f
C457 distortionUnit_3.tgate_1.CTRLB VGND 4.8561f
C458 a_9642_28858# VGND 0.674093f
C459 a_6912_30102# VGND 5.69112f
C460 a_8014_30557# VGND 1.73604f
C461 distortionUnit_3.myOpamp_0.INn VGND 8.10346f
C462 distortionUnit_3.tgate_1.IN VGND 2.63329f
C463 a_7756_30557# VGND 3.01493f
C464 distortionUnit_5.IN VGND 37.692898f
C465 distortionUnit_4.IN VGND 13.2873f
C466 distortionUnit_2.tgate_1.CTRLB VGND 4.829f
C467 a_22410_34902# VGND 0.675619f
C468 a_19680_36146# VGND 5.66142f
C469 a_20782_36601# VGND 1.72068f
C470 distortionUnit_2.myOpamp_0.INn VGND 8.00351f
C471 distortionUnit_2.tgate_1.IN VGND 2.61296f
C472 a_20524_36601# VGND 2.92111f
C473 distortionUnit_1.tgate_1.CTRLB VGND 4.89426f
C474 a_9596_34746# VGND 0.67333f
C475 a_6866_35990# VGND 5.75062f
C476 a_7968_36445# VGND 1.77546f
C477 distortionUnit_1.myOpamp_0.INn VGND 8.23525f
C478 distortionUnit_1.tgate_1.IN VGND 2.71686f
C479 a_7710_36445# VGND 3.45573f
C480 distortionUnit_3.IN VGND 29.620098f
C481 distortionUnit_2.IN VGND 13.223f
C482 distortionUnit_7.sky130_fd_sc_hd__tap_2_0.VPB VGND 1.14309f
C483 distortionUnit_0.sky130_fd_sc_hd__tap_2_0.VPB VGND 1.14329f
C484 distortionUnit_6.sky130_fd_sc_hd__tap_2_0.VPB VGND 1.14329f
C485 distortionUnit_5.sky130_fd_sc_hd__tap_2_0.VPB VGND 1.14329f
C486 distortionUnit_4.sky130_fd_sc_hd__tap_2_0.VPB VGND 1.14329f
C487 distortionUnit_3.sky130_fd_sc_hd__tap_2_0.VPB VGND 1.14329f
C488 distortionUnit_2.sky130_fd_sc_hd__tap_2_0.VPB VGND 1.14329f
C489 distortionUnit_1.sky130_fd_sc_hd__tap_2_0.VPB VGND 1.14329f
C490 ui_in[0].t1 VGND 0.009827f
C491 ui_in[0].t10 VGND 0.005791f
C492 ui_in[0].t6 VGND 0.009827f
C493 ui_in[0].t15 VGND 0.005791f
C494 ui_in[0].n0 VGND 0.014172f
C495 ui_in[0].t3 VGND 0.009827f
C496 ui_in[0].t11 VGND 0.005791f
C497 ui_in[0].t8 VGND 0.009827f
C498 ui_in[0].t16 VGND 0.005791f
C499 ui_in[0].n1 VGND 0.014172f
C500 ui_in[0].t13 VGND 0.009827f
C501 ui_in[0].t18 VGND 0.005791f
C502 ui_in[0].n2 VGND 0.013246f
C503 ui_in[0].n3 VGND 0.006486f
C504 ui_in[0].n4 VGND 0.005382f
C505 ui_in[0].n5 VGND 0.006486f
C506 ui_in[0].n6 VGND 0.014172f
C507 ui_in[0].n7 VGND 0.006486f
C508 ui_in[0].n8 VGND 0.005382f
C509 ui_in[0].n9 VGND 0.005382f
C510 ui_in[0].n10 VGND 0.006486f
C511 ui_in[0].n11 VGND 0.014172f
C512 ui_in[0].t12 VGND 0.009827f
C513 ui_in[0].t17 VGND 0.005791f
C514 ui_in[0].t5 VGND 0.009827f
C515 ui_in[0].t14 VGND 0.005791f
C516 ui_in[0].n12 VGND 0.014172f
C517 ui_in[0].t0 VGND 0.009827f
C518 ui_in[0].t9 VGND 0.005791f
C519 ui_in[0].n13 VGND 0.013246f
C520 ui_in[0].n14 VGND 0.00693f
C521 ui_in[0].n15 VGND 0.005382f
C522 ui_in[0].n16 VGND 0.006486f
C523 ui_in[0].n17 VGND 0.014172f
C524 ui_in[0].n18 VGND 0.006486f
C525 ui_in[0].n19 VGND 0.004855f
C526 ui_in[0].n20 VGND 0.330015f
C527 ui_in[0].t7 VGND 0.106933f
C528 ui_in[0].t2 VGND 0.106932f
C529 ui_in[0].n21 VGND 0.618901f
C530 ui_in[0].n22 VGND 0.406141f
C531 ui_in[0].n23 VGND 2.15842f
C532 ui_in[0].t4 VGND 0.109802f
C533 ui_in[0].t19 VGND 0.109801f
C534 ui_in[0].n24 VGND 0.605904f
C535 ui_in[0].n25 VGND 0.410629f
C536 ui_in[0].n26 VGND 1.14138f
C537 ui_in[1].t10 VGND 0.012664f
C538 ui_in[1].t1 VGND 0.007463f
C539 ui_in[1].t4 VGND 0.012664f
C540 ui_in[1].t12 VGND 0.007463f
C541 ui_in[1].n0 VGND 0.018264f
C542 ui_in[1].t7 VGND 0.012664f
C543 ui_in[1].t17 VGND 0.007463f
C544 ui_in[1].t11 VGND 0.012664f
C545 ui_in[1].t2 VGND 0.007463f
C546 ui_in[1].n1 VGND 0.018264f
C547 ui_in[1].t8 VGND 0.012664f
C548 ui_in[1].t18 VGND 0.007463f
C549 ui_in[1].n2 VGND 0.01707f
C550 ui_in[1].n3 VGND 0.008358f
C551 ui_in[1].n4 VGND 0.006935f
C552 ui_in[1].n5 VGND 0.008358f
C553 ui_in[1].n6 VGND 0.018264f
C554 ui_in[1].n7 VGND 0.008358f
C555 ui_in[1].n8 VGND 0.006935f
C556 ui_in[1].n9 VGND 0.006935f
C557 ui_in[1].n10 VGND 0.008358f
C558 ui_in[1].n11 VGND 0.018264f
C559 ui_in[1].t6 VGND 0.012664f
C560 ui_in[1].t16 VGND 0.007463f
C561 ui_in[1].t9 VGND 0.012664f
C562 ui_in[1].t19 VGND 0.007463f
C563 ui_in[1].n12 VGND 0.018264f
C564 ui_in[1].t5 VGND 0.012664f
C565 ui_in[1].t13 VGND 0.007463f
C566 ui_in[1].n13 VGND 0.01707f
C567 ui_in[1].n14 VGND 0.00893f
C568 ui_in[1].n15 VGND 0.006935f
C569 ui_in[1].n16 VGND 0.008358f
C570 ui_in[1].n17 VGND 0.018264f
C571 ui_in[1].n18 VGND 0.008358f
C572 ui_in[1].n19 VGND 0.006257f
C573 ui_in[1].n20 VGND 0.42528f
C574 ui_in[1].t14 VGND 0.137801f
C575 ui_in[1].t15 VGND 0.137799f
C576 ui_in[1].n21 VGND 0.797557f
C577 ui_in[1].n22 VGND 0.523381f
C578 ui_in[1].n23 VGND 2.78149f
C579 ui_in[1].t0 VGND 0.141499f
C580 ui_in[1].t3 VGND 0.141497f
C581 ui_in[1].n24 VGND 0.780809f
C582 ui_in[1].n25 VGND 0.529164f
C583 ui_in[1].n26 VGND 1.47086f
C584 ui_in[5].t16 VGND 0.012772f
C585 ui_in[5].t7 VGND 0.007526f
C586 ui_in[5].t14 VGND 0.012772f
C587 ui_in[5].t5 VGND 0.007526f
C588 ui_in[5].n0 VGND 0.018418f
C589 ui_in[5].t18 VGND 0.012772f
C590 ui_in[5].t8 VGND 0.007526f
C591 ui_in[5].t0 VGND 0.012772f
C592 ui_in[5].t10 VGND 0.007526f
C593 ui_in[5].n1 VGND 0.018418f
C594 ui_in[5].t19 VGND 0.012772f
C595 ui_in[5].t9 VGND 0.007526f
C596 ui_in[5].n2 VGND 0.017214f
C597 ui_in[5].n3 VGND 0.008429f
C598 ui_in[5].n4 VGND 0.006994f
C599 ui_in[5].n5 VGND 0.008429f
C600 ui_in[5].n6 VGND 0.018418f
C601 ui_in[5].n7 VGND 0.008429f
C602 ui_in[5].n8 VGND 0.006994f
C603 ui_in[5].n9 VGND 0.006994f
C604 ui_in[5].n10 VGND 0.008429f
C605 ui_in[5].n11 VGND 0.018418f
C606 ui_in[5].t11 VGND 0.012772f
C607 ui_in[5].t2 VGND 0.007526f
C608 ui_in[5].t12 VGND 0.012772f
C609 ui_in[5].t3 VGND 0.007526f
C610 ui_in[5].n12 VGND 0.018418f
C611 ui_in[5].t15 VGND 0.012772f
C612 ui_in[5].t6 VGND 0.007526f
C613 ui_in[5].n13 VGND 0.017214f
C614 ui_in[5].n14 VGND 0.009006f
C615 ui_in[5].n15 VGND 0.006994f
C616 ui_in[5].n16 VGND 0.008429f
C617 ui_in[5].n17 VGND 0.018418f
C618 ui_in[5].n18 VGND 0.008429f
C619 ui_in[5].n19 VGND 0.00631f
C620 ui_in[5].n20 VGND 0.428882f
C621 ui_in[5].t4 VGND 0.138968f
C622 ui_in[5].t1 VGND 0.138967f
C623 ui_in[5].n21 VGND 0.804313f
C624 ui_in[5].n22 VGND 0.527814f
C625 ui_in[5].n23 VGND 2.80505f
C626 ui_in[5].t17 VGND 0.142697f
C627 ui_in[5].t13 VGND 0.142695f
C628 ui_in[5].n24 VGND 0.787423f
C629 ui_in[5].n25 VGND 0.533646f
C630 ui_in[5].n26 VGND 1.48332f
C631 ui_in[2].t9 VGND 0.011838f
C632 ui_in[2].t15 VGND 0.006976f
C633 ui_in[2].t4 VGND 0.011838f
C634 ui_in[2].t12 VGND 0.006976f
C635 ui_in[2].n0 VGND 0.017073f
C636 ui_in[2].t10 VGND 0.011838f
C637 ui_in[2].t16 VGND 0.006976f
C638 ui_in[2].t1 VGND 0.011838f
C639 ui_in[2].t7 VGND 0.006976f
C640 ui_in[2].n1 VGND 0.017073f
C641 ui_in[2].t5 VGND 0.011838f
C642 ui_in[2].t13 VGND 0.006976f
C643 ui_in[2].n2 VGND 0.015957f
C644 ui_in[2].n3 VGND 0.007813f
C645 ui_in[2].n4 VGND 0.006483f
C646 ui_in[2].n5 VGND 0.007813f
C647 ui_in[2].n6 VGND 0.017073f
C648 ui_in[2].n7 VGND 0.007813f
C649 ui_in[2].n8 VGND 0.006483f
C650 ui_in[2].n9 VGND 0.006483f
C651 ui_in[2].n10 VGND 0.007813f
C652 ui_in[2].n11 VGND 0.017073f
C653 ui_in[2].t3 VGND 0.011838f
C654 ui_in[2].t11 VGND 0.006976f
C655 ui_in[2].t0 VGND 0.011838f
C656 ui_in[2].t6 VGND 0.006976f
C657 ui_in[2].n12 VGND 0.017073f
C658 ui_in[2].t2 VGND 0.011838f
C659 ui_in[2].t8 VGND 0.006976f
C660 ui_in[2].n13 VGND 0.015957f
C661 ui_in[2].n14 VGND 0.008348f
C662 ui_in[2].n15 VGND 0.006483f
C663 ui_in[2].n16 VGND 0.007813f
C664 ui_in[2].n17 VGND 0.017073f
C665 ui_in[2].n18 VGND 0.007813f
C666 ui_in[2].n19 VGND 0.005849f
C667 ui_in[2].n20 VGND 0.39755f
C668 ui_in[2].t18 VGND 0.128816f
C669 ui_in[2].t19 VGND 0.128814f
C670 ui_in[2].n21 VGND 0.745554f
C671 ui_in[2].n22 VGND 0.489254f
C672 ui_in[2].n23 VGND 2.60012f
C673 ui_in[2].t14 VGND 0.132272f
C674 ui_in[2].t17 VGND 0.132271f
C675 ui_in[2].n24 VGND 0.729898f
C676 ui_in[2].n25 VGND 0.494661f
C677 ui_in[2].n26 VGND 1.37496f
C678 ua[0].t4 VGND 0.044597f
C679 ua[0].t8 VGND 0.04445f
C680 ua[0].n0 VGND 0.055058f
C681 ua[0].t6 VGND 0.04445f
C682 ua[0].n1 VGND 0.032483f
C683 ua[0].t5 VGND 0.04445f
C684 ua[0].n2 VGND 0.028193f
C685 ua[0].t7 VGND 0.044564f
C686 ua[0].n3 VGND 0.077301f
C687 ua[0].t0 VGND 0.010208f
C688 ua[0].n4 VGND 0.039441f
C689 ua[0].t2 VGND 0.002822f
C690 ua[0].t3 VGND 0.002822f
C691 ua[0].n5 VGND 0.009159f
C692 ua[0].n6 VGND 0.055852f
C693 ua[0].t1 VGND 0.010208f
C694 ua[0].n7 VGND 0.029466f
C695 ua[0].n8 VGND 0.33763f
C696 ua[0].n9 VGND 0.814452f
C697 ua[0].n10 VGND 0.409633f
C698 ua[0].n11 VGND 0.158424f
C699 ua[1].n0 VGND 0.043178f
C700 ua[1].t3 VGND 0.001064f
C701 ua[1].t2 VGND 0.001064f
C702 ua[1].n1 VGND 0.002204f
C703 ua[1].t6 VGND 0.003846f
C704 ua[1].n2 VGND 0.030935f
C705 ua[1].n3 VGND 0.028972f
C706 ua[1].t7 VGND 0.003805f
C707 ua[1].n4 VGND 0.030242f
C708 ua[1].n5 VGND 0.097005f
C709 ua[1].n6 VGND 0.043178f
C710 ua[1].t4 VGND 0.001064f
C711 ua[1].t5 VGND 0.001064f
C712 ua[1].n7 VGND 0.002204f
C713 ua[1].t0 VGND 0.003846f
C714 ua[1].n8 VGND 0.030935f
C715 ua[1].n9 VGND 0.028972f
C716 ua[1].t1 VGND 0.003805f
C717 ua[1].n10 VGND 0.030242f
C718 ua[1].n11 VGND 0.075781f
C719 ua[1].n12 VGND 0.199199f
C720 ua[1].n13 VGND 1.7979f
C721 ui_in[7].t8 VGND 0.010065f
C722 ui_in[7].t17 VGND 0.005931f
C723 ui_in[7].t4 VGND 0.010065f
C724 ui_in[7].t14 VGND 0.005931f
C725 ui_in[7].n0 VGND 0.014515f
C726 ui_in[7].t3 VGND 0.010065f
C727 ui_in[7].t13 VGND 0.005931f
C728 ui_in[7].t9 VGND 0.010065f
C729 ui_in[7].t18 VGND 0.005931f
C730 ui_in[7].n1 VGND 0.014515f
C731 ui_in[7].t5 VGND 0.010065f
C732 ui_in[7].t15 VGND 0.005931f
C733 ui_in[7].n2 VGND 0.013566f
C734 ui_in[7].n3 VGND 0.006643f
C735 ui_in[7].n4 VGND 0.005512f
C736 ui_in[7].n5 VGND 0.006643f
C737 ui_in[7].n6 VGND 0.014515f
C738 ui_in[7].n7 VGND 0.006643f
C739 ui_in[7].n8 VGND 0.005512f
C740 ui_in[7].n9 VGND 0.005512f
C741 ui_in[7].n10 VGND 0.006643f
C742 ui_in[7].n11 VGND 0.014515f
C743 ui_in[7].t2 VGND 0.010065f
C744 ui_in[7].t12 VGND 0.005931f
C745 ui_in[7].t6 VGND 0.010065f
C746 ui_in[7].t16 VGND 0.005931f
C747 ui_in[7].n12 VGND 0.014515f
C748 ui_in[7].t1 VGND 0.010065f
C749 ui_in[7].t11 VGND 0.005931f
C750 ui_in[7].n13 VGND 0.013566f
C751 ui_in[7].n14 VGND 0.007098f
C752 ui_in[7].n15 VGND 0.005512f
C753 ui_in[7].n16 VGND 0.006643f
C754 ui_in[7].n17 VGND 0.014515f
C755 ui_in[7].n18 VGND 0.006643f
C756 ui_in[7].n19 VGND 0.004973f
C757 ui_in[7].n20 VGND 0.337994f
C758 ui_in[7].t7 VGND 0.109518f
C759 ui_in[7].t10 VGND 0.109517f
C760 ui_in[7].n21 VGND 0.633864f
C761 ui_in[7].n22 VGND 0.41596f
C762 ui_in[7].n23 VGND 2.2106f
C763 ui_in[7].t19 VGND 0.112457f
C764 ui_in[7].t0 VGND 0.112455f
C765 ui_in[7].n24 VGND 0.620553f
C766 ui_in[7].n25 VGND 0.420556f
C767 ui_in[7].n26 VGND 1.16898f
C768 distortionUnit_5.IN.t14 VGND 0.04871f
C769 distortionUnit_5.IN.t13 VGND 0.048551f
C770 distortionUnit_5.IN.n0 VGND 0.060137f
C771 distortionUnit_5.IN.t15 VGND 0.048551f
C772 distortionUnit_5.IN.n1 VGND 0.03548f
C773 distortionUnit_5.IN.t16 VGND 0.048551f
C774 distortionUnit_5.IN.n2 VGND 0.030794f
C775 distortionUnit_5.IN.t12 VGND 0.048675f
C776 distortionUnit_5.IN.n3 VGND 0.084432f
C777 distortionUnit_5.IN.t4 VGND 0.011149f
C778 distortionUnit_5.IN.n4 VGND 0.04308f
C779 distortionUnit_5.IN.t10 VGND 0.003083f
C780 distortionUnit_5.IN.t11 VGND 0.003083f
C781 distortionUnit_5.IN.n5 VGND 0.010004f
C782 distortionUnit_5.IN.n6 VGND 0.061004f
C783 distortionUnit_5.IN.t5 VGND 0.011149f
C784 distortionUnit_5.IN.n7 VGND 0.032184f
C785 distortionUnit_5.IN.n8 VGND 0.368775f
C786 distortionUnit_5.IN.n9 VGND 1.41753f
C787 distortionUnit_5.IN.n10 VGND 5.86744f
C788 distortionUnit_5.IN.n11 VGND 0.125118f
C789 distortionUnit_5.IN.t7 VGND 0.003083f
C790 distortionUnit_5.IN.t6 VGND 0.003083f
C791 distortionUnit_5.IN.n12 VGND 0.006386f
C792 distortionUnit_5.IN.t1 VGND 0.011144f
C793 distortionUnit_5.IN.n13 VGND 0.089641f
C794 distortionUnit_5.IN.n14 VGND 0.083951f
C795 distortionUnit_5.IN.t0 VGND 0.011026f
C796 distortionUnit_5.IN.n15 VGND 0.087633f
C797 distortionUnit_5.IN.n16 VGND 0.281094f
C798 distortionUnit_5.IN.n17 VGND 0.577223f
C799 distortionUnit_5.IN.n18 VGND 0.219593f
C800 distortionUnit_5.IN.t9 VGND 0.011026f
C801 distortionUnit_5.IN.n19 VGND 0.087633f
C802 distortionUnit_5.IN.t3 VGND 0.003083f
C803 distortionUnit_5.IN.t2 VGND 0.003083f
C804 distortionUnit_5.IN.n20 VGND 0.006386f
C805 distortionUnit_5.IN.n21 VGND 0.083951f
C806 distortionUnit_5.IN.t8 VGND 0.011144f
C807 distortionUnit_5.IN.n22 VGND 0.089641f
C808 distortionUnit_5.IN.n23 VGND 0.125118f
C809 ui_in[3].t8 VGND 0.01219f
C810 ui_in[3].t18 VGND 0.007184f
C811 ui_in[3].t12 VGND 0.01219f
C812 ui_in[3].t2 VGND 0.007184f
C813 ui_in[3].n0 VGND 0.01758f
C814 ui_in[3].t16 VGND 0.01219f
C815 ui_in[3].t6 VGND 0.007184f
C816 ui_in[3].t15 VGND 0.01219f
C817 ui_in[3].t5 VGND 0.007184f
C818 ui_in[3].n1 VGND 0.01758f
C819 ui_in[3].t17 VGND 0.01219f
C820 ui_in[3].t7 VGND 0.007184f
C821 ui_in[3].n2 VGND 0.016431f
C822 ui_in[3].n3 VGND 0.008046f
C823 ui_in[3].n4 VGND 0.006676f
C824 ui_in[3].n5 VGND 0.008046f
C825 ui_in[3].n6 VGND 0.01758f
C826 ui_in[3].n7 VGND 0.008046f
C827 ui_in[3].n8 VGND 0.006676f
C828 ui_in[3].n9 VGND 0.006676f
C829 ui_in[3].n10 VGND 0.008046f
C830 ui_in[3].n11 VGND 0.01758f
C831 ui_in[3].t9 VGND 0.01219f
C832 ui_in[3].t19 VGND 0.007184f
C833 ui_in[3].t11 VGND 0.01219f
C834 ui_in[3].t1 VGND 0.007184f
C835 ui_in[3].n12 VGND 0.01758f
C836 ui_in[3].t13 VGND 0.01219f
C837 ui_in[3].t3 VGND 0.007184f
C838 ui_in[3].n13 VGND 0.016431f
C839 ui_in[3].n14 VGND 0.008596f
C840 ui_in[3].n15 VGND 0.006676f
C841 ui_in[3].n16 VGND 0.008046f
C842 ui_in[3].n17 VGND 0.01758f
C843 ui_in[3].n18 VGND 0.008046f
C844 ui_in[3].n19 VGND 0.006023f
C845 ui_in[3].n20 VGND 0.409367f
C846 ui_in[3].t14 VGND 0.132645f
C847 ui_in[3].t4 VGND 0.132643f
C848 ui_in[3].n21 VGND 0.767714f
C849 ui_in[3].n22 VGND 0.503797f
C850 ui_in[3].n23 VGND 2.67741f
C851 ui_in[3].t0 VGND 0.136204f
C852 ui_in[3].t10 VGND 0.136202f
C853 ui_in[3].n24 VGND 0.751592f
C854 ui_in[3].n25 VGND 0.509363f
C855 ui_in[3].n26 VGND 1.41582f
C856 ui_in[6].t5 VGND 0.013589f
C857 ui_in[6].t15 VGND 0.008008f
C858 ui_in[6].t7 VGND 0.013589f
C859 ui_in[6].t17 VGND 0.008008f
C860 ui_in[6].n0 VGND 0.019597f
C861 ui_in[6].t6 VGND 0.013589f
C862 ui_in[6].t16 VGND 0.008008f
C863 ui_in[6].t4 VGND 0.013589f
C864 ui_in[6].t14 VGND 0.008008f
C865 ui_in[6].n1 VGND 0.019597f
C866 ui_in[6].t1 VGND 0.013589f
C867 ui_in[6].t12 VGND 0.008008f
C868 ui_in[6].n2 VGND 0.018316f
C869 ui_in[6].n3 VGND 0.008969f
C870 ui_in[6].n4 VGND 0.007442f
C871 ui_in[6].n5 VGND 0.008969f
C872 ui_in[6].n6 VGND 0.019597f
C873 ui_in[6].n7 VGND 0.008969f
C874 ui_in[6].n8 VGND 0.007442f
C875 ui_in[6].n9 VGND 0.007442f
C876 ui_in[6].n10 VGND 0.008969f
C877 ui_in[6].n11 VGND 0.019597f
C878 ui_in[6].t0 VGND 0.013589f
C879 ui_in[6].t11 VGND 0.008008f
C880 ui_in[6].t2 VGND 0.013589f
C881 ui_in[6].t13 VGND 0.008008f
C882 ui_in[6].n12 VGND 0.019597f
C883 ui_in[6].t18 VGND 0.013589f
C884 ui_in[6].t9 VGND 0.008008f
C885 ui_in[6].n13 VGND 0.018316f
C886 ui_in[6].n14 VGND 0.009583f
C887 ui_in[6].n15 VGND 0.007442f
C888 ui_in[6].n16 VGND 0.008969f
C889 ui_in[6].n17 VGND 0.019597f
C890 ui_in[6].n18 VGND 0.008969f
C891 ui_in[6].n19 VGND 0.006714f
C892 ui_in[6].n20 VGND 0.456338f
C893 ui_in[6].t8 VGND 0.147865f
C894 ui_in[6].t10 VGND 0.147863f
C895 ui_in[6].n21 VGND 0.855802f
C896 ui_in[6].n22 VGND 0.561603f
C897 ui_in[6].n23 VGND 2.98462f
C898 ui_in[6].t19 VGND 0.151832f
C899 ui_in[6].t3 VGND 0.15183f
C900 ui_in[6].n24 VGND 0.837831f
C901 ui_in[6].n25 VGND 0.567808f
C902 ui_in[6].n26 VGND 1.57828f
C903 VPWR.n0 VGND 0.623237f
C904 VPWR.n1 VGND 0.674759f
C905 VPWR.n2 VGND 0.110507f
C906 VPWR.n3 VGND 0.110453f
C907 VPWR.n4 VGND 0.221041f
C908 VPWR.n5 VGND 0.221205f
C909 VPWR.n6 VGND 0.671834f
C910 VPWR.n7 VGND 0.110398f
C911 VPWR.n8 VGND 0.110753f
C912 VPWR.n9 VGND 0.66017f
C913 VPWR.n10 VGND 0.110104f
C914 VPWR.n11 VGND 0.109753f
C915 VPWR.n12 VGND 0.21972f
C916 VPWR.n13 VGND 0.659318f
C917 VPWR.n14 VGND 0.674341f
C918 VPWR.n15 VGND 0.661022f
C919 VPWR.n16 VGND 0.21994f
C920 VPWR.n17 VGND 0.109942f
C921 VPWR.n18 VGND 0.109996f
C922 VPWR.n19 VGND 0.378218f
C923 VPWR.n20 VGND 0.705663f
C924 VPWR.t259 VGND 0.038722f
C925 VPWR.t261 VGND 0.008769f
C926 VPWR.n21 VGND 0.050741f
C927 VPWR.t210 VGND 0.002387f
C928 VPWR.t194 VGND 0.002387f
C929 VPWR.n22 VGND 0.004935f
C930 VPWR.n23 VGND 0.098003f
C931 VPWR.t198 VGND 0.002387f
C932 VPWR.t202 VGND 0.002387f
C933 VPWR.n24 VGND 0.004935f
C934 VPWR.n25 VGND 0.082388f
C935 VPWR.t250 VGND 0.038696f
C936 VPWR.t252 VGND 0.008769f
C937 VPWR.n26 VGND 0.090592f
C938 VPWR.t200 VGND 0.002387f
C939 VPWR.t204 VGND 0.002387f
C940 VPWR.n27 VGND 0.004935f
C941 VPWR.n28 VGND 0.119479f
C942 VPWR.t212 VGND 0.002387f
C943 VPWR.t196 VGND 0.002387f
C944 VPWR.n29 VGND 0.004935f
C945 VPWR.n30 VGND 0.072018f
C946 VPWR.t260 VGND 0.136104f
C947 VPWR.t209 VGND 0.108715f
C948 VPWR.t193 VGND 0.108715f
C949 VPWR.t197 VGND 0.108715f
C950 VPWR.t201 VGND 0.108715f
C951 VPWR.t207 VGND 0.078165f
C952 VPWR.t251 VGND 0.136104f
C953 VPWR.t203 VGND 0.108715f
C954 VPWR.t199 VGND 0.108715f
C955 VPWR.t195 VGND 0.108715f
C956 VPWR.t211 VGND 0.108715f
C957 VPWR.t205 VGND 0.084907f
C958 VPWR.n31 VGND -0.063754f
C959 VPWR.t3 VGND 0.091568f
C960 VPWR.n32 VGND 0.14066f
C961 VPWR.n33 VGND 0.018764f
C962 VPWR.t208 VGND 0.002387f
C963 VPWR.t206 VGND 0.002387f
C964 VPWR.n34 VGND 0.004935f
C965 VPWR.n35 VGND 0.08098f
C966 VPWR.n36 VGND 2.88464f
C967 VPWR.n37 VGND 1.41734f
C968 VPWR.n38 VGND 0.003792f
C969 VPWR.n39 VGND 0.007269f
C970 VPWR.t84 VGND 0.002222f
C971 VPWR.t79 VGND 0.002222f
C972 VPWR.n40 VGND 0.00477f
C973 VPWR.t305 VGND 0.002222f
C974 VPWR.t87 VGND 0.002222f
C975 VPWR.n41 VGND 0.00477f
C976 VPWR.n42 VGND 0.001987f
C977 VPWR.t82 VGND 0.00846f
C978 VPWR.n43 VGND 0.012053f
C979 VPWR.n44 VGND 0.005452f
C980 VPWR.n45 VGND 0.007269f
C981 VPWR.n46 VGND 0.007269f
C982 VPWR.n47 VGND 0.001413f
C983 VPWR.n48 VGND 0.005438f
C984 VPWR.n49 VGND 0.00235f
C985 VPWR.n50 VGND 0.005438f
C986 VPWR.t136 VGND 0.002222f
C987 VPWR.t20 VGND 0.002222f
C988 VPWR.n51 VGND 0.00477f
C989 VPWR.n52 VGND 0.001791f
C990 VPWR.t192 VGND 0.008461f
C991 VPWR.n53 VGND 0.009943f
C992 VPWR.n54 VGND 0.004534f
C993 VPWR.n55 VGND 0.007269f
C994 VPWR.n56 VGND 0.007269f
C995 VPWR.n57 VGND 0.001609f
C996 VPWR.n58 VGND 0.005438f
C997 VPWR.n59 VGND 0.002253f
C998 VPWR.n60 VGND 0.001385f
C999 VPWR.n61 VGND 0.007111f
C1000 VPWR.n62 VGND 0.292138f
C1001 VPWR.n63 VGND 0.029053f
C1002 VPWR.n64 VGND 0.016745f
C1003 VPWR.n65 VGND 0.119512f
C1004 VPWR.t25 VGND 0.095282f
C1005 VPWR.n66 VGND 0.060303f
C1006 VPWR.t184 VGND 0.095282f
C1007 VPWR.n67 VGND 0.098727f
C1008 VPWR.n68 VGND 0.051668f
C1009 VPWR.n69 VGND 0.227646f
C1010 VPWR.n70 VGND 0.029053f
C1011 VPWR.n71 VGND 0.016745f
C1012 VPWR.n72 VGND 0.119512f
C1013 VPWR.t131 VGND 0.095282f
C1014 VPWR.n73 VGND 0.060303f
C1015 VPWR.t132 VGND 0.095282f
C1016 VPWR.n74 VGND 0.098727f
C1017 VPWR.n75 VGND 0.051668f
C1018 VPWR.n76 VGND 0.230467f
C1019 VPWR.n77 VGND 0.212137f
C1020 VPWR.n78 VGND 29.499098f
C1021 VPWR.n79 VGND 0.623237f
C1022 VPWR.n80 VGND 0.674759f
C1023 VPWR.n81 VGND 0.110507f
C1024 VPWR.n82 VGND 0.110453f
C1025 VPWR.n83 VGND 0.221041f
C1026 VPWR.n84 VGND 0.221205f
C1027 VPWR.n85 VGND 0.671834f
C1028 VPWR.n86 VGND 0.110398f
C1029 VPWR.n87 VGND 0.110753f
C1030 VPWR.n88 VGND 0.66017f
C1031 VPWR.n89 VGND 0.110104f
C1032 VPWR.n90 VGND 0.109753f
C1033 VPWR.n91 VGND 0.21972f
C1034 VPWR.n92 VGND 0.659318f
C1035 VPWR.n93 VGND 0.674341f
C1036 VPWR.n94 VGND 0.661022f
C1037 VPWR.n95 VGND 0.21994f
C1038 VPWR.n96 VGND 0.109942f
C1039 VPWR.n97 VGND 0.109996f
C1040 VPWR.n98 VGND 0.378218f
C1041 VPWR.n99 VGND 0.705663f
C1042 VPWR.t247 VGND 0.038722f
C1043 VPWR.t249 VGND 0.008769f
C1044 VPWR.n100 VGND 0.050741f
C1045 VPWR.t93 VGND 0.002387f
C1046 VPWR.t95 VGND 0.002387f
C1047 VPWR.n101 VGND 0.004935f
C1048 VPWR.n102 VGND 0.098003f
C1049 VPWR.t103 VGND 0.002387f
C1050 VPWR.t101 VGND 0.002387f
C1051 VPWR.n103 VGND 0.004935f
C1052 VPWR.n104 VGND 0.082388f
C1053 VPWR.t256 VGND 0.038696f
C1054 VPWR.t258 VGND 0.008769f
C1055 VPWR.n105 VGND 0.090592f
C1056 VPWR.t97 VGND 0.002387f
C1057 VPWR.t105 VGND 0.002387f
C1058 VPWR.n106 VGND 0.004935f
C1059 VPWR.n107 VGND 0.119479f
C1060 VPWR.t91 VGND 0.002387f
C1061 VPWR.t99 VGND 0.002387f
C1062 VPWR.n108 VGND 0.004935f
C1063 VPWR.n109 VGND 0.072018f
C1064 VPWR.t248 VGND 0.136104f
C1065 VPWR.t92 VGND 0.108715f
C1066 VPWR.t94 VGND 0.108715f
C1067 VPWR.t102 VGND 0.108715f
C1068 VPWR.t100 VGND 0.108715f
C1069 VPWR.t106 VGND 0.078165f
C1070 VPWR.t257 VGND 0.136104f
C1071 VPWR.t104 VGND 0.108715f
C1072 VPWR.t96 VGND 0.108715f
C1073 VPWR.t98 VGND 0.108715f
C1074 VPWR.t90 VGND 0.108715f
C1075 VPWR.t108 VGND 0.084907f
C1076 VPWR.n110 VGND -0.063754f
C1077 VPWR.t187 VGND 0.091568f
C1078 VPWR.n111 VGND 0.14066f
C1079 VPWR.n112 VGND 0.018764f
C1080 VPWR.t107 VGND 0.002387f
C1081 VPWR.t109 VGND 0.002387f
C1082 VPWR.n113 VGND 0.004935f
C1083 VPWR.n114 VGND 0.08098f
C1084 VPWR.n115 VGND 2.88464f
C1085 VPWR.n116 VGND 1.41734f
C1086 VPWR.n117 VGND 0.003792f
C1087 VPWR.n118 VGND 0.007269f
C1088 VPWR.t159 VGND 0.002222f
C1089 VPWR.t80 VGND 0.002222f
C1090 VPWR.n119 VGND 0.00477f
C1091 VPWR.t52 VGND 0.002222f
C1092 VPWR.t54 VGND 0.002222f
C1093 VPWR.n120 VGND 0.00477f
C1094 VPWR.n121 VGND 0.001987f
C1095 VPWR.t306 VGND 0.00846f
C1096 VPWR.n122 VGND 0.012053f
C1097 VPWR.n123 VGND 0.005452f
C1098 VPWR.n124 VGND 0.007269f
C1099 VPWR.n125 VGND 0.007269f
C1100 VPWR.n126 VGND 0.001413f
C1101 VPWR.n127 VGND 0.005438f
C1102 VPWR.n128 VGND 0.00235f
C1103 VPWR.n129 VGND 0.005438f
C1104 VPWR.t21 VGND 0.002222f
C1105 VPWR.t5 VGND 0.002222f
C1106 VPWR.n130 VGND 0.00477f
C1107 VPWR.n131 VGND 0.001791f
C1108 VPWR.t307 VGND 0.008461f
C1109 VPWR.n132 VGND 0.009943f
C1110 VPWR.n133 VGND 0.004534f
C1111 VPWR.n134 VGND 0.007269f
C1112 VPWR.n135 VGND 0.007269f
C1113 VPWR.n136 VGND 0.001609f
C1114 VPWR.n137 VGND 0.005438f
C1115 VPWR.n138 VGND 0.002253f
C1116 VPWR.n139 VGND 0.001385f
C1117 VPWR.n140 VGND 0.007111f
C1118 VPWR.n141 VGND 0.292138f
C1119 VPWR.n142 VGND 0.029053f
C1120 VPWR.n143 VGND 0.016745f
C1121 VPWR.n144 VGND 0.119512f
C1122 VPWR.t88 VGND 0.095282f
C1123 VPWR.n145 VGND 0.060303f
C1124 VPWR.t86 VGND 0.095282f
C1125 VPWR.n146 VGND 0.098727f
C1126 VPWR.n147 VGND 0.051668f
C1127 VPWR.n148 VGND 0.227646f
C1128 VPWR.n149 VGND 0.029053f
C1129 VPWR.n150 VGND 0.016745f
C1130 VPWR.n151 VGND 0.119512f
C1131 VPWR.t181 VGND 0.095282f
C1132 VPWR.n152 VGND 0.060303f
C1133 VPWR.t180 VGND 0.095282f
C1134 VPWR.n153 VGND 0.098727f
C1135 VPWR.n154 VGND 0.051668f
C1136 VPWR.n155 VGND 0.230467f
C1137 VPWR.n156 VGND 0.212137f
C1138 VPWR.n157 VGND 5.02724f
C1139 VPWR.n158 VGND 0.414202p
C1140 VPWR.n159 VGND 15.4034f
C1141 VPWR.n160 VGND 0.623237f
C1142 VPWR.n161 VGND 0.674759f
C1143 VPWR.n162 VGND 0.110507f
C1144 VPWR.n163 VGND 0.110453f
C1145 VPWR.n164 VGND 0.221041f
C1146 VPWR.n165 VGND 0.221205f
C1147 VPWR.n166 VGND 0.671834f
C1148 VPWR.n167 VGND 0.110398f
C1149 VPWR.n168 VGND 0.110753f
C1150 VPWR.n169 VGND 0.66017f
C1151 VPWR.n170 VGND 0.110104f
C1152 VPWR.n171 VGND 0.109753f
C1153 VPWR.n172 VGND 0.21972f
C1154 VPWR.n173 VGND 0.659318f
C1155 VPWR.n174 VGND 0.674341f
C1156 VPWR.n175 VGND 0.661022f
C1157 VPWR.n176 VGND 0.21994f
C1158 VPWR.n177 VGND 0.109942f
C1159 VPWR.n178 VGND 0.109996f
C1160 VPWR.n179 VGND 0.378218f
C1161 VPWR.n180 VGND 0.705663f
C1162 VPWR.t241 VGND 0.038722f
C1163 VPWR.t243 VGND 0.008769f
C1164 VPWR.n181 VGND 0.050741f
C1165 VPWR.t144 VGND 0.002387f
C1166 VPWR.t150 VGND 0.002387f
C1167 VPWR.n182 VGND 0.004935f
C1168 VPWR.n183 VGND 0.098003f
C1169 VPWR.t154 VGND 0.002387f
C1170 VPWR.t142 VGND 0.002387f
C1171 VPWR.n184 VGND 0.004935f
C1172 VPWR.n185 VGND 0.082388f
C1173 VPWR.t238 VGND 0.038696f
C1174 VPWR.t240 VGND 0.008769f
C1175 VPWR.n186 VGND 0.090592f
C1176 VPWR.t138 VGND 0.002387f
C1177 VPWR.t156 VGND 0.002387f
C1178 VPWR.n187 VGND 0.004935f
C1179 VPWR.n188 VGND 0.119479f
C1180 VPWR.t148 VGND 0.002387f
C1181 VPWR.t152 VGND 0.002387f
C1182 VPWR.n189 VGND 0.004935f
C1183 VPWR.n190 VGND 0.072018f
C1184 VPWR.t242 VGND 0.136104f
C1185 VPWR.t143 VGND 0.108715f
C1186 VPWR.t149 VGND 0.108715f
C1187 VPWR.t153 VGND 0.108715f
C1188 VPWR.t141 VGND 0.108715f
C1189 VPWR.t139 VGND 0.078165f
C1190 VPWR.t239 VGND 0.136104f
C1191 VPWR.t155 VGND 0.108715f
C1192 VPWR.t137 VGND 0.108715f
C1193 VPWR.t151 VGND 0.108715f
C1194 VPWR.t147 VGND 0.108715f
C1195 VPWR.t145 VGND 0.084907f
C1196 VPWR.n191 VGND -0.063754f
C1197 VPWR.t83 VGND 0.091568f
C1198 VPWR.n192 VGND 0.14066f
C1199 VPWR.n193 VGND 0.018764f
C1200 VPWR.t140 VGND 0.002387f
C1201 VPWR.t146 VGND 0.002387f
C1202 VPWR.n194 VGND 0.004935f
C1203 VPWR.n195 VGND 0.08098f
C1204 VPWR.n196 VGND 2.88464f
C1205 VPWR.n197 VGND 1.41734f
C1206 VPWR.n198 VGND 0.003792f
C1207 VPWR.n199 VGND 0.007269f
C1208 VPWR.t303 VGND 0.002222f
C1209 VPWR.t0 VGND 0.002222f
C1210 VPWR.n200 VGND 0.00477f
C1211 VPWR.t12 VGND 0.002222f
C1212 VPWR.t85 VGND 0.002222f
C1213 VPWR.n201 VGND 0.00477f
C1214 VPWR.n202 VGND 0.001987f
C1215 VPWR.t27 VGND 0.00846f
C1216 VPWR.n203 VGND 0.012053f
C1217 VPWR.n204 VGND 0.005452f
C1218 VPWR.n205 VGND 0.007269f
C1219 VPWR.n206 VGND 0.007269f
C1220 VPWR.n207 VGND 0.001413f
C1221 VPWR.n208 VGND 0.005438f
C1222 VPWR.n209 VGND 0.00235f
C1223 VPWR.n210 VGND 0.005438f
C1224 VPWR.t53 VGND 0.002222f
C1225 VPWR.t89 VGND 0.002222f
C1226 VPWR.n211 VGND 0.00477f
C1227 VPWR.n212 VGND 0.001791f
C1228 VPWR.t1 VGND 0.008461f
C1229 VPWR.n213 VGND 0.009943f
C1230 VPWR.n214 VGND 0.004534f
C1231 VPWR.n215 VGND 0.007269f
C1232 VPWR.n216 VGND 0.007269f
C1233 VPWR.n217 VGND 0.001609f
C1234 VPWR.n218 VGND 0.005438f
C1235 VPWR.n219 VGND 0.002253f
C1236 VPWR.n220 VGND 0.001385f
C1237 VPWR.n221 VGND 0.007111f
C1238 VPWR.n222 VGND 0.292138f
C1239 VPWR.n223 VGND 0.029053f
C1240 VPWR.n224 VGND 0.016745f
C1241 VPWR.n225 VGND 0.119512f
C1242 VPWR.t189 VGND 0.095282f
C1243 VPWR.n226 VGND 0.060303f
C1244 VPWR.t190 VGND 0.095282f
C1245 VPWR.n227 VGND 0.098727f
C1246 VPWR.n228 VGND 0.051668f
C1247 VPWR.n229 VGND 0.227646f
C1248 VPWR.n230 VGND 0.029053f
C1249 VPWR.n231 VGND 0.016745f
C1250 VPWR.n232 VGND 0.119512f
C1251 VPWR.t28 VGND 0.095282f
C1252 VPWR.n233 VGND 0.060303f
C1253 VPWR.t29 VGND 0.095282f
C1254 VPWR.n234 VGND 0.098727f
C1255 VPWR.n235 VGND 0.051668f
C1256 VPWR.n236 VGND 0.230467f
C1257 VPWR.n237 VGND 0.212137f
C1258 VPWR.n238 VGND 12.623199f
C1259 VPWR.n239 VGND 0.623237f
C1260 VPWR.n240 VGND 0.674759f
C1261 VPWR.n241 VGND 0.110507f
C1262 VPWR.n242 VGND 0.110453f
C1263 VPWR.n243 VGND 0.221041f
C1264 VPWR.n244 VGND 0.221205f
C1265 VPWR.n245 VGND 0.671834f
C1266 VPWR.n246 VGND 0.110398f
C1267 VPWR.n247 VGND 0.110753f
C1268 VPWR.n248 VGND 0.66017f
C1269 VPWR.n249 VGND 0.110104f
C1270 VPWR.n250 VGND 0.109753f
C1271 VPWR.n251 VGND 0.21972f
C1272 VPWR.n252 VGND 0.659318f
C1273 VPWR.n253 VGND 0.674341f
C1274 VPWR.n254 VGND 0.661022f
C1275 VPWR.n255 VGND 0.21994f
C1276 VPWR.n256 VGND 0.109942f
C1277 VPWR.n257 VGND 0.109996f
C1278 VPWR.n258 VGND 0.378218f
C1279 VPWR.n259 VGND 0.705663f
C1280 VPWR.t229 VGND 0.038722f
C1281 VPWR.t231 VGND 0.008769f
C1282 VPWR.n260 VGND 0.050741f
C1283 VPWR.t165 VGND 0.002387f
C1284 VPWR.t169 VGND 0.002387f
C1285 VPWR.n261 VGND 0.004935f
C1286 VPWR.n262 VGND 0.098003f
C1287 VPWR.t175 VGND 0.002387f
C1288 VPWR.t161 VGND 0.002387f
C1289 VPWR.n263 VGND 0.004935f
C1290 VPWR.n264 VGND 0.082388f
C1291 VPWR.t235 VGND 0.038696f
C1292 VPWR.t237 VGND 0.008769f
C1293 VPWR.n265 VGND 0.090592f
C1294 VPWR.t171 VGND 0.002387f
C1295 VPWR.t177 VGND 0.002387f
C1296 VPWR.n266 VGND 0.004935f
C1297 VPWR.n267 VGND 0.119479f
C1298 VPWR.t167 VGND 0.002387f
C1299 VPWR.t173 VGND 0.002387f
C1300 VPWR.n268 VGND 0.004935f
C1301 VPWR.n269 VGND 0.072018f
C1302 VPWR.t230 VGND 0.136104f
C1303 VPWR.t164 VGND 0.108715f
C1304 VPWR.t168 VGND 0.108715f
C1305 VPWR.t174 VGND 0.108715f
C1306 VPWR.t160 VGND 0.108715f
C1307 VPWR.t178 VGND 0.078165f
C1308 VPWR.t236 VGND 0.136104f
C1309 VPWR.t176 VGND 0.108715f
C1310 VPWR.t170 VGND 0.108715f
C1311 VPWR.t172 VGND 0.108715f
C1312 VPWR.t166 VGND 0.108715f
C1313 VPWR.t162 VGND 0.084907f
C1314 VPWR.n270 VGND -0.063754f
C1315 VPWR.t26 VGND 0.091568f
C1316 VPWR.n271 VGND 0.14066f
C1317 VPWR.n272 VGND 0.018764f
C1318 VPWR.t179 VGND 0.002387f
C1319 VPWR.t163 VGND 0.002387f
C1320 VPWR.n273 VGND 0.004935f
C1321 VPWR.n274 VGND 0.08098f
C1322 VPWR.n275 VGND 2.88464f
C1323 VPWR.n276 VGND 1.41734f
C1324 VPWR.n277 VGND 0.003792f
C1325 VPWR.n278 VGND 0.007269f
C1326 VPWR.t188 VGND 0.002222f
C1327 VPWR.t14 VGND 0.002222f
C1328 VPWR.n279 VGND 0.00477f
C1329 VPWR.t274 VGND 0.002222f
C1330 VPWR.t298 VGND 0.002222f
C1331 VPWR.n280 VGND 0.00477f
C1332 VPWR.n281 VGND 0.001987f
C1333 VPWR.t301 VGND 0.00846f
C1334 VPWR.n282 VGND 0.012053f
C1335 VPWR.n283 VGND 0.005452f
C1336 VPWR.n284 VGND 0.007269f
C1337 VPWR.n285 VGND 0.007269f
C1338 VPWR.n286 VGND 0.001413f
C1339 VPWR.n287 VGND 0.005438f
C1340 VPWR.n288 VGND 0.00235f
C1341 VPWR.n289 VGND 0.005438f
C1342 VPWR.t275 VGND 0.002222f
C1343 VPWR.t81 VGND 0.002222f
C1344 VPWR.n290 VGND 0.00477f
C1345 VPWR.n291 VGND 0.001791f
C1346 VPWR.t130 VGND 0.008461f
C1347 VPWR.n292 VGND 0.009943f
C1348 VPWR.n293 VGND 0.004534f
C1349 VPWR.n294 VGND 0.007269f
C1350 VPWR.n295 VGND 0.007269f
C1351 VPWR.n296 VGND 0.001609f
C1352 VPWR.n297 VGND 0.005438f
C1353 VPWR.n298 VGND 0.002253f
C1354 VPWR.n299 VGND 0.001385f
C1355 VPWR.n300 VGND 0.007111f
C1356 VPWR.n301 VGND 0.292138f
C1357 VPWR.n302 VGND 0.029053f
C1358 VPWR.n303 VGND 0.016745f
C1359 VPWR.n304 VGND 0.119512f
C1360 VPWR.t6 VGND 0.095282f
C1361 VPWR.n305 VGND 0.060303f
C1362 VPWR.t133 VGND 0.095282f
C1363 VPWR.n306 VGND 0.098727f
C1364 VPWR.n307 VGND 0.051668f
C1365 VPWR.n308 VGND 0.227646f
C1366 VPWR.n309 VGND 0.029053f
C1367 VPWR.n310 VGND 0.016745f
C1368 VPWR.n311 VGND 0.119512f
C1369 VPWR.t308 VGND 0.095282f
C1370 VPWR.n312 VGND 0.060303f
C1371 VPWR.t309 VGND 0.095282f
C1372 VPWR.n313 VGND 0.098727f
C1373 VPWR.n314 VGND 0.051668f
C1374 VPWR.n315 VGND 0.230467f
C1375 VPWR.n316 VGND 0.212137f
C1376 VPWR.n317 VGND 5.02724f
C1377 VPWR.n318 VGND 0.346099p
C1378 VPWR.n319 VGND 0.029053f
C1379 VPWR.n320 VGND 0.016745f
C1380 VPWR.n321 VGND 0.119512f
C1381 VPWR.t77 VGND 0.095282f
C1382 VPWR.n322 VGND 0.060303f
C1383 VPWR.t76 VGND 0.095282f
C1384 VPWR.n323 VGND 0.098727f
C1385 VPWR.n324 VGND 0.051668f
C1386 VPWR.n325 VGND 0.227646f
C1387 VPWR.n326 VGND 0.029053f
C1388 VPWR.n327 VGND 0.016745f
C1389 VPWR.n328 VGND 0.119512f
C1390 VPWR.t272 VGND 0.095282f
C1391 VPWR.n329 VGND 0.060303f
C1392 VPWR.t273 VGND 0.095282f
C1393 VPWR.n330 VGND 0.098727f
C1394 VPWR.n331 VGND 0.051668f
C1395 VPWR.n332 VGND 0.230467f
C1396 VPWR.n333 VGND 0.511231f
C1397 VPWR.n334 VGND 0.003792f
C1398 VPWR.n335 VGND 0.007269f
C1399 VPWR.t135 VGND 0.002222f
C1400 VPWR.t18 VGND 0.002222f
C1401 VPWR.n336 VGND 0.00477f
C1402 VPWR.t78 VGND 0.002222f
C1403 VPWR.t304 VGND 0.002222f
C1404 VPWR.n337 VGND 0.00477f
C1405 VPWR.n338 VGND 0.001987f
C1406 VPWR.t51 VGND 0.00846f
C1407 VPWR.n339 VGND 0.012053f
C1408 VPWR.n340 VGND 0.005452f
C1409 VPWR.n341 VGND 0.007269f
C1410 VPWR.n342 VGND 0.007269f
C1411 VPWR.n343 VGND 0.001413f
C1412 VPWR.n344 VGND 0.005438f
C1413 VPWR.n345 VGND 0.00235f
C1414 VPWR.n346 VGND 0.005438f
C1415 VPWR.t75 VGND 0.002222f
C1416 VPWR.t19 VGND 0.002222f
C1417 VPWR.n347 VGND 0.00477f
C1418 VPWR.n348 VGND 0.001791f
C1419 VPWR.t15 VGND 0.008461f
C1420 VPWR.n349 VGND 0.009943f
C1421 VPWR.n350 VGND 0.004534f
C1422 VPWR.n351 VGND 0.007269f
C1423 VPWR.n352 VGND 0.007269f
C1424 VPWR.n353 VGND 0.001609f
C1425 VPWR.n354 VGND 0.005438f
C1426 VPWR.n355 VGND 0.002253f
C1427 VPWR.n356 VGND 0.001385f
C1428 VPWR.n357 VGND 0.007111f
C1429 VPWR.n358 VGND 0.292138f
C1430 VPWR.n359 VGND 7.26512f
C1431 VPWR.n360 VGND 0.623237f
C1432 VPWR.n361 VGND 0.674759f
C1433 VPWR.n362 VGND 0.110507f
C1434 VPWR.n363 VGND 0.110453f
C1435 VPWR.n364 VGND 0.221041f
C1436 VPWR.n365 VGND 0.221205f
C1437 VPWR.n366 VGND 0.671834f
C1438 VPWR.n367 VGND 0.110398f
C1439 VPWR.n368 VGND 0.110753f
C1440 VPWR.n369 VGND 0.66017f
C1441 VPWR.n370 VGND 0.110104f
C1442 VPWR.n371 VGND 0.109753f
C1443 VPWR.n372 VGND 0.21972f
C1444 VPWR.n373 VGND 0.659318f
C1445 VPWR.n374 VGND 0.674341f
C1446 VPWR.n375 VGND 0.661022f
C1447 VPWR.n376 VGND 0.21994f
C1448 VPWR.n377 VGND 0.109942f
C1449 VPWR.n378 VGND 0.109996f
C1450 VPWR.n379 VGND 0.378218f
C1451 VPWR.n380 VGND 0.705663f
C1452 VPWR.t226 VGND 0.038722f
C1453 VPWR.t228 VGND 0.008769f
C1454 VPWR.n381 VGND 0.050741f
C1455 VPWR.t286 VGND 0.002387f
C1456 VPWR.t284 VGND 0.002387f
C1457 VPWR.n382 VGND 0.004935f
C1458 VPWR.n383 VGND 0.098003f
C1459 VPWR.t290 VGND 0.002387f
C1460 VPWR.t278 VGND 0.002387f
C1461 VPWR.n384 VGND 0.004935f
C1462 VPWR.n385 VGND 0.082388f
C1463 VPWR.t232 VGND 0.038696f
C1464 VPWR.t234 VGND 0.008769f
C1465 VPWR.n386 VGND 0.090592f
C1466 VPWR.t292 VGND 0.002387f
C1467 VPWR.t294 VGND 0.002387f
C1468 VPWR.n387 VGND 0.004935f
C1469 VPWR.n388 VGND 0.119479f
C1470 VPWR.t280 VGND 0.002387f
C1471 VPWR.t288 VGND 0.002387f
C1472 VPWR.n389 VGND 0.004935f
C1473 VPWR.n390 VGND 0.072018f
C1474 VPWR.t227 VGND 0.136104f
C1475 VPWR.t285 VGND 0.108715f
C1476 VPWR.t283 VGND 0.108715f
C1477 VPWR.t289 VGND 0.108715f
C1478 VPWR.t277 VGND 0.108715f
C1479 VPWR.t295 VGND 0.078165f
C1480 VPWR.t233 VGND 0.136104f
C1481 VPWR.t293 VGND 0.108715f
C1482 VPWR.t291 VGND 0.108715f
C1483 VPWR.t287 VGND 0.108715f
C1484 VPWR.t279 VGND 0.108715f
C1485 VPWR.t281 VGND 0.084907f
C1486 VPWR.n391 VGND -0.063754f
C1487 VPWR.t186 VGND 0.091568f
C1488 VPWR.n392 VGND 0.14066f
C1489 VPWR.n393 VGND 0.018764f
C1490 VPWR.t296 VGND 0.002387f
C1491 VPWR.t282 VGND 0.002387f
C1492 VPWR.n394 VGND 0.004935f
C1493 VPWR.n395 VGND 0.08098f
C1494 VPWR.n396 VGND 2.88464f
C1495 VPWR.n397 VGND 1.41734f
C1496 VPWR.n398 VGND 4.93141f
C1497 VPWR.n399 VGND 0.029053f
C1498 VPWR.n400 VGND 0.016745f
C1499 VPWR.n401 VGND 0.119512f
C1500 VPWR.t221 VGND 0.095282f
C1501 VPWR.n402 VGND 0.060303f
C1502 VPWR.t213 VGND 0.095282f
C1503 VPWR.n403 VGND 0.098727f
C1504 VPWR.n404 VGND 0.051668f
C1505 VPWR.n405 VGND 0.227646f
C1506 VPWR.n406 VGND 0.029053f
C1507 VPWR.n407 VGND 0.016745f
C1508 VPWR.n408 VGND 0.119512f
C1509 VPWR.t311 VGND 0.095282f
C1510 VPWR.n409 VGND 0.060303f
C1511 VPWR.t310 VGND 0.095282f
C1512 VPWR.n410 VGND 0.098727f
C1513 VPWR.n411 VGND 0.051668f
C1514 VPWR.n412 VGND 0.230467f
C1515 VPWR.n413 VGND 0.212137f
C1516 VPWR.n414 VGND 3.43552f
C1517 VPWR.n415 VGND 0.003792f
C1518 VPWR.n416 VGND 0.007269f
C1519 VPWR.t219 VGND 0.002222f
C1520 VPWR.t217 VGND 0.002222f
C1521 VPWR.n417 VGND 0.00477f
C1522 VPWR.t216 VGND 0.002222f
C1523 VPWR.t214 VGND 0.002222f
C1524 VPWR.n418 VGND 0.00477f
C1525 VPWR.n419 VGND 0.001987f
C1526 VPWR.t218 VGND 0.00846f
C1527 VPWR.n420 VGND 0.012053f
C1528 VPWR.n421 VGND 0.005452f
C1529 VPWR.n422 VGND 0.007269f
C1530 VPWR.n423 VGND 0.007269f
C1531 VPWR.n424 VGND 0.001413f
C1532 VPWR.n425 VGND 0.005438f
C1533 VPWR.n426 VGND 0.00235f
C1534 VPWR.n427 VGND 0.005438f
C1535 VPWR.t220 VGND 0.002222f
C1536 VPWR.t222 VGND 0.002222f
C1537 VPWR.n428 VGND 0.00477f
C1538 VPWR.n429 VGND 0.001791f
C1539 VPWR.t215 VGND 0.008461f
C1540 VPWR.n430 VGND 0.009943f
C1541 VPWR.n431 VGND 0.004534f
C1542 VPWR.n432 VGND 0.007269f
C1543 VPWR.n433 VGND 0.007269f
C1544 VPWR.n434 VGND 0.001609f
C1545 VPWR.n435 VGND 0.005438f
C1546 VPWR.n436 VGND 0.002253f
C1547 VPWR.n437 VGND 0.001385f
C1548 VPWR.n438 VGND 0.007111f
C1549 VPWR.n439 VGND 0.292138f
C1550 VPWR.n440 VGND 4.83713f
C1551 VPWR.n441 VGND 0.623237f
C1552 VPWR.n442 VGND 0.674759f
C1553 VPWR.n443 VGND 0.110507f
C1554 VPWR.n444 VGND 0.110453f
C1555 VPWR.n445 VGND 0.221041f
C1556 VPWR.n446 VGND 0.221205f
C1557 VPWR.n447 VGND 0.671834f
C1558 VPWR.n448 VGND 0.110398f
C1559 VPWR.n449 VGND 0.110753f
C1560 VPWR.n450 VGND 0.66017f
C1561 VPWR.n451 VGND 0.110104f
C1562 VPWR.n452 VGND 0.109753f
C1563 VPWR.n453 VGND 0.21972f
C1564 VPWR.n454 VGND 0.659318f
C1565 VPWR.n455 VGND 0.674341f
C1566 VPWR.n456 VGND 0.661022f
C1567 VPWR.n457 VGND 0.21994f
C1568 VPWR.n458 VGND 0.109942f
C1569 VPWR.n459 VGND 0.109996f
C1570 VPWR.n460 VGND 0.378218f
C1571 VPWR.n461 VGND 0.705663f
C1572 VPWR.t223 VGND 0.038722f
C1573 VPWR.t225 VGND 0.008769f
C1574 VPWR.n462 VGND 0.050741f
C1575 VPWR.t66 VGND 0.002387f
C1576 VPWR.t70 VGND 0.002387f
C1577 VPWR.n463 VGND 0.004935f
C1578 VPWR.n464 VGND 0.098003f
C1579 VPWR.t74 VGND 0.002387f
C1580 VPWR.t62 VGND 0.002387f
C1581 VPWR.n465 VGND 0.004935f
C1582 VPWR.n466 VGND 0.082388f
C1583 VPWR.t244 VGND 0.038696f
C1584 VPWR.t246 VGND 0.008769f
C1585 VPWR.n467 VGND 0.090592f
C1586 VPWR.t58 VGND 0.002387f
C1587 VPWR.t56 VGND 0.002387f
C1588 VPWR.n468 VGND 0.004935f
C1589 VPWR.n469 VGND 0.119479f
C1590 VPWR.t64 VGND 0.002387f
C1591 VPWR.t72 VGND 0.002387f
C1592 VPWR.n470 VGND 0.004935f
C1593 VPWR.n471 VGND 0.072018f
C1594 VPWR.t224 VGND 0.136104f
C1595 VPWR.t65 VGND 0.108715f
C1596 VPWR.t69 VGND 0.108715f
C1597 VPWR.t73 VGND 0.108715f
C1598 VPWR.t61 VGND 0.108715f
C1599 VPWR.t59 VGND 0.078165f
C1600 VPWR.t245 VGND 0.136104f
C1601 VPWR.t55 VGND 0.108715f
C1602 VPWR.t57 VGND 0.108715f
C1603 VPWR.t71 VGND 0.108715f
C1604 VPWR.t63 VGND 0.108715f
C1605 VPWR.t67 VGND 0.084907f
C1606 VPWR.n472 VGND -0.063754f
C1607 VPWR.t182 VGND 0.091568f
C1608 VPWR.n473 VGND 0.14066f
C1609 VPWR.n474 VGND 0.018764f
C1610 VPWR.t60 VGND 0.002387f
C1611 VPWR.t68 VGND 0.002387f
C1612 VPWR.n475 VGND 0.004935f
C1613 VPWR.n476 VGND 0.08098f
C1614 VPWR.n477 VGND 2.88464f
C1615 VPWR.n478 VGND 1.41734f
C1616 VPWR.n479 VGND 4.93141f
C1617 VPWR.n480 VGND 7.56566f
C1618 VPWR.n481 VGND 0.029053f
C1619 VPWR.n482 VGND 0.016745f
C1620 VPWR.n483 VGND 0.119512f
C1621 VPWR.t17 VGND 0.095282f
C1622 VPWR.n484 VGND 0.060303f
C1623 VPWR.t134 VGND 0.095282f
C1624 VPWR.n485 VGND 0.098727f
C1625 VPWR.n486 VGND 0.051668f
C1626 VPWR.n487 VGND 0.227646f
C1627 VPWR.n488 VGND 0.029053f
C1628 VPWR.n489 VGND 0.016745f
C1629 VPWR.n490 VGND 0.119512f
C1630 VPWR.t157 VGND 0.095282f
C1631 VPWR.n491 VGND 0.060303f
C1632 VPWR.t158 VGND 0.095282f
C1633 VPWR.n492 VGND 0.098727f
C1634 VPWR.n493 VGND 0.051668f
C1635 VPWR.n494 VGND 0.230467f
C1636 VPWR.n495 VGND 0.451918f
C1637 VPWR.n496 VGND 0.003792f
C1638 VPWR.n497 VGND 0.007269f
C1639 VPWR.t16 VGND 0.002222f
C1640 VPWR.t302 VGND 0.002222f
C1641 VPWR.n498 VGND 0.00477f
C1642 VPWR.t299 VGND 0.002222f
C1643 VPWR.t191 VGND 0.002222f
C1644 VPWR.n499 VGND 0.00477f
C1645 VPWR.n500 VGND 0.001987f
C1646 VPWR.t50 VGND 0.00846f
C1647 VPWR.n501 VGND 0.012053f
C1648 VPWR.n502 VGND 0.005452f
C1649 VPWR.n503 VGND 0.007269f
C1650 VPWR.n504 VGND 0.007269f
C1651 VPWR.n505 VGND 0.001413f
C1652 VPWR.n506 VGND 0.005438f
C1653 VPWR.n507 VGND 0.00235f
C1654 VPWR.n508 VGND 0.005438f
C1655 VPWR.t300 VGND 0.002222f
C1656 VPWR.t7 VGND 0.002222f
C1657 VPWR.n509 VGND 0.00477f
C1658 VPWR.n510 VGND 0.001791f
C1659 VPWR.t24 VGND 0.008461f
C1660 VPWR.n511 VGND 0.009943f
C1661 VPWR.n512 VGND 0.004534f
C1662 VPWR.n513 VGND 0.007269f
C1663 VPWR.n514 VGND 0.007269f
C1664 VPWR.n515 VGND 0.001609f
C1665 VPWR.n516 VGND 0.005438f
C1666 VPWR.n517 VGND 0.002253f
C1667 VPWR.n518 VGND 0.001385f
C1668 VPWR.n519 VGND 0.007111f
C1669 VPWR.n520 VGND 0.292138f
C1670 VPWR.n521 VGND 5.28636f
C1671 VPWR.n522 VGND 0.623237f
C1672 VPWR.n523 VGND 0.674759f
C1673 VPWR.n524 VGND 0.110507f
C1674 VPWR.n525 VGND 0.110453f
C1675 VPWR.n526 VGND 0.221041f
C1676 VPWR.n527 VGND 0.221205f
C1677 VPWR.n528 VGND 0.671834f
C1678 VPWR.n529 VGND 0.110398f
C1679 VPWR.n530 VGND 0.110753f
C1680 VPWR.n531 VGND 0.66017f
C1681 VPWR.n532 VGND 0.110104f
C1682 VPWR.n533 VGND 0.109753f
C1683 VPWR.n534 VGND 0.21972f
C1684 VPWR.n535 VGND 0.659318f
C1685 VPWR.n536 VGND 0.674341f
C1686 VPWR.n537 VGND 0.661022f
C1687 VPWR.n538 VGND 0.21994f
C1688 VPWR.n539 VGND 0.109942f
C1689 VPWR.n540 VGND 0.109996f
C1690 VPWR.n541 VGND 0.378218f
C1691 VPWR.n542 VGND 0.705663f
C1692 VPWR.t262 VGND 0.038722f
C1693 VPWR.t264 VGND 0.008769f
C1694 VPWR.n543 VGND 0.050741f
C1695 VPWR.t127 VGND 0.002387f
C1696 VPWR.t113 VGND 0.002387f
C1697 VPWR.n544 VGND 0.004935f
C1698 VPWR.n545 VGND 0.098003f
C1699 VPWR.t115 VGND 0.002387f
C1700 VPWR.t119 VGND 0.002387f
C1701 VPWR.n546 VGND 0.004935f
C1702 VPWR.n547 VGND 0.082388f
C1703 VPWR.t253 VGND 0.038696f
C1704 VPWR.t255 VGND 0.008769f
C1705 VPWR.n548 VGND 0.090592f
C1706 VPWR.t117 VGND 0.002387f
C1707 VPWR.t121 VGND 0.002387f
C1708 VPWR.n549 VGND 0.004935f
C1709 VPWR.n550 VGND 0.119479f
C1710 VPWR.t111 VGND 0.002387f
C1711 VPWR.t129 VGND 0.002387f
C1712 VPWR.n551 VGND 0.004935f
C1713 VPWR.n552 VGND 0.072018f
C1714 VPWR.t263 VGND 0.136104f
C1715 VPWR.t126 VGND 0.108715f
C1716 VPWR.t112 VGND 0.108715f
C1717 VPWR.t114 VGND 0.108715f
C1718 VPWR.t118 VGND 0.108715f
C1719 VPWR.t124 VGND 0.078165f
C1720 VPWR.t254 VGND 0.136104f
C1721 VPWR.t120 VGND 0.108715f
C1722 VPWR.t116 VGND 0.108715f
C1723 VPWR.t128 VGND 0.108715f
C1724 VPWR.t110 VGND 0.108715f
C1725 VPWR.t122 VGND 0.084907f
C1726 VPWR.n553 VGND -0.063754f
C1727 VPWR.t13 VGND 0.091568f
C1728 VPWR.n554 VGND 0.14066f
C1729 VPWR.n555 VGND 0.018764f
C1730 VPWR.t125 VGND 0.002387f
C1731 VPWR.t123 VGND 0.002387f
C1732 VPWR.n556 VGND 0.004935f
C1733 VPWR.n557 VGND 0.08098f
C1734 VPWR.n558 VGND 2.88464f
C1735 VPWR.n559 VGND 1.41734f
C1736 VPWR.n560 VGND 3.69855f
C1737 VPWR.n561 VGND 0.029053f
C1738 VPWR.n562 VGND 0.016745f
C1739 VPWR.n563 VGND 0.119512f
C1740 VPWR.t4 VGND 0.095282f
C1741 VPWR.n564 VGND 0.060303f
C1742 VPWR.t22 VGND 0.095282f
C1743 VPWR.n565 VGND 0.098727f
C1744 VPWR.n566 VGND 0.051668f
C1745 VPWR.n567 VGND 0.227646f
C1746 VPWR.n568 VGND 0.029053f
C1747 VPWR.n569 VGND 0.016745f
C1748 VPWR.n570 VGND 0.119512f
C1749 VPWR.t8 VGND 0.095282f
C1750 VPWR.n571 VGND 0.060303f
C1751 VPWR.t9 VGND 0.095282f
C1752 VPWR.n572 VGND 0.098727f
C1753 VPWR.n573 VGND 0.051668f
C1754 VPWR.n574 VGND 0.230467f
C1755 VPWR.n575 VGND 0.212137f
C1756 VPWR.n576 VGND 2.8107f
C1757 VPWR.n577 VGND 0.003792f
C1758 VPWR.n578 VGND 0.007269f
C1759 VPWR.t23 VGND 0.002222f
C1760 VPWR.t297 VGND 0.002222f
C1761 VPWR.n579 VGND 0.00477f
C1762 VPWR.t10 VGND 0.002222f
C1763 VPWR.t11 VGND 0.002222f
C1764 VPWR.n580 VGND 0.00477f
C1765 VPWR.n581 VGND 0.001987f
C1766 VPWR.t185 VGND 0.00846f
C1767 VPWR.n582 VGND 0.012053f
C1768 VPWR.n583 VGND 0.005452f
C1769 VPWR.n584 VGND 0.007269f
C1770 VPWR.n585 VGND 0.007269f
C1771 VPWR.n586 VGND 0.001413f
C1772 VPWR.n587 VGND 0.005438f
C1773 VPWR.n588 VGND 0.00235f
C1774 VPWR.n589 VGND 0.005438f
C1775 VPWR.t271 VGND 0.002222f
C1776 VPWR.t2 VGND 0.002222f
C1777 VPWR.n590 VGND 0.00477f
C1778 VPWR.n591 VGND 0.001791f
C1779 VPWR.t183 VGND 0.008461f
C1780 VPWR.n592 VGND 0.009943f
C1781 VPWR.n593 VGND 0.004534f
C1782 VPWR.n594 VGND 0.007269f
C1783 VPWR.n595 VGND 0.007269f
C1784 VPWR.n596 VGND 0.001609f
C1785 VPWR.n597 VGND 0.005438f
C1786 VPWR.n598 VGND 0.002253f
C1787 VPWR.n599 VGND 0.001385f
C1788 VPWR.n600 VGND 0.007111f
C1789 VPWR.n601 VGND 0.292138f
C1790 VPWR.n602 VGND 3.82649f
C1791 VPWR.n603 VGND 0.623237f
C1792 VPWR.n604 VGND 0.674759f
C1793 VPWR.n605 VGND 0.110507f
C1794 VPWR.n606 VGND 0.110453f
C1795 VPWR.n607 VGND 0.221041f
C1796 VPWR.n608 VGND 0.221205f
C1797 VPWR.n609 VGND 0.671834f
C1798 VPWR.n610 VGND 0.110398f
C1799 VPWR.n611 VGND 0.110753f
C1800 VPWR.n612 VGND 0.66017f
C1801 VPWR.n613 VGND 0.110104f
C1802 VPWR.n614 VGND 0.109753f
C1803 VPWR.n615 VGND 0.21972f
C1804 VPWR.n616 VGND 0.659318f
C1805 VPWR.n617 VGND 0.674341f
C1806 VPWR.n618 VGND 0.661022f
C1807 VPWR.n619 VGND 0.21994f
C1808 VPWR.n620 VGND 0.109942f
C1809 VPWR.n621 VGND 0.109996f
C1810 VPWR.n622 VGND 0.378218f
C1811 VPWR.n623 VGND 0.705663f
C1812 VPWR.t268 VGND 0.038722f
C1813 VPWR.t270 VGND 0.008769f
C1814 VPWR.n624 VGND 0.050741f
C1815 VPWR.t47 VGND 0.002387f
C1816 VPWR.t37 VGND 0.002387f
C1817 VPWR.n625 VGND 0.004935f
C1818 VPWR.n626 VGND 0.098003f
C1819 VPWR.t35 VGND 0.002387f
C1820 VPWR.t41 VGND 0.002387f
C1821 VPWR.n627 VGND 0.004935f
C1822 VPWR.n628 VGND 0.082388f
C1823 VPWR.t265 VGND 0.038696f
C1824 VPWR.t267 VGND 0.008769f
C1825 VPWR.n629 VGND 0.090592f
C1826 VPWR.t39 VGND 0.002387f
C1827 VPWR.t43 VGND 0.002387f
C1828 VPWR.n630 VGND 0.004935f
C1829 VPWR.n631 VGND 0.119479f
C1830 VPWR.t33 VGND 0.002387f
C1831 VPWR.t31 VGND 0.002387f
C1832 VPWR.n632 VGND 0.004935f
C1833 VPWR.n633 VGND 0.072018f
C1834 VPWR.t269 VGND 0.136104f
C1835 VPWR.t46 VGND 0.108715f
C1836 VPWR.t36 VGND 0.108715f
C1837 VPWR.t34 VGND 0.108715f
C1838 VPWR.t40 VGND 0.108715f
C1839 VPWR.t44 VGND 0.078165f
C1840 VPWR.t266 VGND 0.136104f
C1841 VPWR.t42 VGND 0.108715f
C1842 VPWR.t38 VGND 0.108715f
C1843 VPWR.t30 VGND 0.108715f
C1844 VPWR.t32 VGND 0.108715f
C1845 VPWR.t48 VGND 0.084907f
C1846 VPWR.n634 VGND -0.063754f
C1847 VPWR.t276 VGND 0.091568f
C1848 VPWR.n635 VGND 0.14066f
C1849 VPWR.n636 VGND 0.018764f
C1850 VPWR.t45 VGND 0.002387f
C1851 VPWR.t49 VGND 0.002387f
C1852 VPWR.n637 VGND 0.004935f
C1853 VPWR.n638 VGND 0.08098f
C1854 VPWR.n639 VGND 2.88464f
C1855 VPWR.n640 VGND 1.41734f
C1856 VPWR.n641 VGND 3.69855f
C1857 VPWR.n642 VGND 7.15614f
C1858 ui_in[4].t10 VGND 0.012697f
C1859 ui_in[4].t0 VGND 0.007482f
C1860 ui_in[4].t8 VGND 0.012697f
C1861 ui_in[4].t18 VGND 0.007482f
C1862 ui_in[4].n0 VGND 0.018311f
C1863 ui_in[4].t15 VGND 0.012697f
C1864 ui_in[4].t4 VGND 0.007482f
C1865 ui_in[4].t13 VGND 0.012697f
C1866 ui_in[4].t2 VGND 0.007482f
C1867 ui_in[4].n1 VGND 0.018311f
C1868 ui_in[4].t9 VGND 0.012697f
C1869 ui_in[4].t19 VGND 0.007482f
C1870 ui_in[4].n2 VGND 0.017114f
C1871 ui_in[4].n3 VGND 0.00838f
C1872 ui_in[4].n4 VGND 0.006953f
C1873 ui_in[4].n5 VGND 0.00838f
C1874 ui_in[4].n6 VGND 0.018311f
C1875 ui_in[4].n7 VGND 0.00838f
C1876 ui_in[4].n8 VGND 0.006953f
C1877 ui_in[4].n9 VGND 0.006953f
C1878 ui_in[4].n10 VGND 0.00838f
C1879 ui_in[4].n11 VGND 0.018311f
C1880 ui_in[4].t7 VGND 0.012697f
C1881 ui_in[4].t17 VGND 0.007482f
C1882 ui_in[4].t5 VGND 0.012697f
C1883 ui_in[4].t11 VGND 0.007482f
C1884 ui_in[4].n12 VGND 0.018311f
C1885 ui_in[4].t14 VGND 0.012697f
C1886 ui_in[4].t3 VGND 0.007482f
C1887 ui_in[4].n13 VGND 0.017114f
C1888 ui_in[4].n14 VGND 0.008954f
C1889 ui_in[4].n15 VGND 0.006953f
C1890 ui_in[4].n16 VGND 0.00838f
C1891 ui_in[4].n17 VGND 0.018311f
C1892 ui_in[4].n18 VGND 0.00838f
C1893 ui_in[4].n19 VGND 0.006273f
C1894 ui_in[4].n20 VGND 0.426388f
C1895 ui_in[4].t1 VGND 0.13816f
C1896 ui_in[4].t12 VGND 0.138158f
C1897 ui_in[4].n21 VGND 0.799636f
C1898 ui_in[4].n22 VGND 0.524745f
C1899 ui_in[4].n23 VGND 2.78873f
C1900 ui_in[4].t16 VGND 0.141867f
C1901 ui_in[4].t6 VGND 0.141865f
C1902 ui_in[4].n24 VGND 0.782844f
C1903 ui_in[4].n25 VGND 0.530543f
C1904 ui_in[4].n26 VGND 1.47469f
.ends

